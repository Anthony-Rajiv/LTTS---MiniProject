dac.sp SPICE FILE
.model nenh nmos
+ level = 2
+   vto = 0.62249   kp = 6.32664e-05   gamma = 0.639243
+   phi = 0.31
+
+   cgso = 2.89e-10   cgdo = 2.89e-10
+   rsh = 60   cj = 0.000327
+   mj = 1.067   cjsw = 1.74e-10   mjsw = 0.195
+   tox = 2.25e-08   nsub = 1.066e+16
+   nss = 3e+10   nfs = 4.55168e+12   tpg = 1
+   xj = 9e-07   ld = 0   uo = 1215.74
+   ucrit = 174667   uexp = 0.0461235
+   vmax = 177269   neff = 4.6883
+
+   delta = 0
.model penh pmos
+ level = 2
+   vto = -0.63025   kp = 2.63544e-05   gamma = 0.618101
+   phi = 0.541111
+
+   cgso = 3.35e-10   cgdo = 3.35e-10
+   rsh = 150   cj = 0.000475
+   mj = 0.341   cjsw = 2.23e-10   mjsw = 0.307
+   tox = 2.25e-08   nsub = 6.57544e+16
+   nss = 3e+10   nfs = 1.66844e+11   tpg = -1
+   xj = 1.12799e-07   ld = 3e-08   uo = 361.941
+   ucrit = 637449   uexp = 0.0888696
+   vmax = 63253.3   neff = 0.64354
+
+   delta = 0
.subckt CMP 1 2 3 4 5
+ 6 7 8 9
md1 10 4 3 9 penh l=5e-07 w=4.8e-06 
+ as=5.27999e-12 ad=2.24e-12 ps=7e-06 pd=3e-06 
+ nrs=0.229167 nrd=0.0972222 
md2 11 5 10 9 penh l=5e-07 w=4.8e-06 
+ as=2.24e-12 ad=4.31999e-12 ps=3e-06 pd=6.6e-06 
+ nrs=0.0972222 nrd=0.1875 
md3 6 8 10 9 penh l=5e-07 w=4.8e-06 
+ as=2.24e-12 ad=4.31999e-12 ps=3e-06 pd=6.6e-06 
+ nrs=0.0972222 nrd=0.1875 
md4 2 11 11 7 nenh l=5e-07 w=2.4e-06 
+ as=1.92e-12 ad=3.84e-12 ps=4.2e-06 pd=5.6e-06 
+ nrs=0.333333 nrd=0.666666 
md5 2 11 6 7 nenh l=5e-07 w=2.4e-06 
+ as=1.92e-12 ad=3.84e-12 ps=4.2e-06 pd=5.6e-06 
+ nrs=0.333333 nrd=0.666666 
c1 2 7 1.14593e-12
c2 6 7 3.3125e-13
c3 7 11 4.02e-13
c4 7 8 6.74875e-13
c5 5 7 2.76104e-13
c6 7 10 8e-18
c7 4 7 4.13662e-13
c8 3 7 1.3488e-12
c9 3 8 1.5e-13
c10 2 10 3.825e-14
c11 2 11 1.4625e-14
c12 5 10 1.4575e-13
c13 6 8 6.6528e-14
c14 5 11 8.175e-14
c15 2 3 3.165e-13
c16 2 8 4.125e-13
c17 3 5 2.955e-13
c18 4 10 1.42e-13
c19 4 11 9e-15
c20 5 8 2e-14
c21 2 6 3.4875e-13
c22 3 4 5.7e-14
c23 4 8 3.5e-14
c24 2 5 4.35e-14
c25 4 6 6.375e-14
c26 3 10 3.825e-14
c27 3 11 2.76375e-13
c28 2 4 2.845e-13
c29 11 8 1.47312e-13
c30 4 5 1.5e-14
.ends CMP
.subckt z2xCMP 1 2 3 4 5
+ 6 7 8 9 10 11
xCMP#1 9 10 2 7 11
+ 6 1 4 2 CMP
xCMP#0 8 10 2 7 11
+ 5 1 3 2 CMP
.ends z2xCMP
.subckt AVddRtg 1 2 3
c31 1 2 6.9264e-12
.ends AVddRtg
.subckt FlashLatchBlnk 1 2 3 4 5
+ 6
c32 1 4 2.9244e-13
c33 1 5 2.69976e-13
c34 1 2 2.68104e-13
c35 1 3 2.88288e-13
c36 5 6 2.1e-14
c37 2 6 2.1e-14
c38 3 6 2.1e-14
c39 4 6 2.1e-14
.ends FlashLatchBlnk
.subckt FlashLatch 1 2 3 4 5
+ 6 7 8 9 10
md6 11 12 10 10 penh l=2e-07 w=2.2e-06 
+ as=1.81396e-12 ad=1.01e-12 ps=3.81886e-06 pd=3.8e-06 
+ nrs=0.374785 nrd=0.208678 
md7 4 13 10 10 penh l=2e-07 w=2.2e-06 
+ as=1.81396e-12 ad=1.01e-12 ps=3.81886e-06 pd=3.8e-06 
+ nrs=0.374785 nrd=0.208678 
md8 14 1 10 10 penh l=2e-07 w=1.8e-06 
+ as=1.48415e-12 ad=7.41598e-13 ps=3.12453e-06 pd=2.23199e-06 
+ nrs=0.458071 nrd=0.228889 
md9 10 11 15 10 penh l=2e-07 w=2.2e-06 
+ as=1.00222e-12 ad=1.81396e-12 ps=3.42221e-06 pd=3.81886e-06 
+ nrs=0.207071 nrd=0.374785 
md10 10 4 3 10 penh l=2e-07 w=2.2e-06 
+ as=8.19309e-13 ad=1.81396e-12 ps=2.50344e-06 pd=3.81886e-06 
+ nrs=0.169279 nrd=0.374785 
md11 11 12 2 2 nenh l=2e-07 w=1.1e-06 
+ as=1.30942e-12 ad=8.79999e-13 ps=4.01923e-06 pd=2.7e-06 
+ nrs=1.08216 nrd=0.727272 
md12 12 5 14 2 nenh l=2e-07 w=7e-07 
+ as=3.40666e-13 ad=3.15e-13 ps=9.79999e-07 pd=9e-07 
+ nrs=0.695237 nrd=0.642857 
md13 15 6 12 2 nenh l=2e-07 w=7e-07 
+ as=3.15e-13 ad=3.66799e-13 ps=9e-07 pd=1.26e-06 
+ nrs=0.642857 nrd=0.74857 
md14 12 6 14 10 penh l=2e-07 w=7e-07 
+ as=2.884e-13 ad=3.15e-13 ps=8.67999e-07 pd=9e-07 
+ nrs=0.588571 nrd=0.642857 
md15 15 5 12 10 penh l=2e-07 w=7e-07 
+ as=3.15e-13 ad=3.18888e-13 ps=9e-07 pd=1.08889e-06 
+ nrs=0.642857 nrd=0.650793 
md16 4 13 2 2 nenh l=2e-07 w=1.1e-06 
+ as=1.30942e-12 ad=8.79999e-13 ps=4.01923e-06 pd=2.7e-06 
+ nrs=1.08216 nrd=0.727272 
md17 13 7 15 2 nenh l=2e-07 w=7e-07 
+ as=3.66799e-13 ad=3.15e-13 ps=1.26e-06 pd=9e-07 
+ nrs=0.74857 nrd=0.642857 
md18 3 8 13 2 nenh l=2e-07 w=7e-07 
+ as=3.15e-13 ad=2.91666e-13 ps=9e-07 pd=8.55554e-07 
+ nrs=0.642857 nrd=0.595238 
md19 13 8 15 10 penh l=2e-07 w=7e-07 
+ as=3.18888e-13 ad=3.15e-13 ps=1.08889e-06 pd=9e-07 
+ nrs=0.650793 nrd=0.642857 
md20 3 7 13 10 penh l=2e-07 w=7e-07 
+ as=3.15e-13 ad=2.60689e-13 ps=9e-07 pd=7.96551e-07 
+ nrs=0.642857 nrd=0.532019 
md21 14 1 2 2 nenh l=2e-07 w=7.99999e-07 
+ as=9.52306e-13 ad=3.89332e-13 ps=2.92307e-06 pd=1.12e-06 
+ nrs=1.48798 nrd=0.608333 
md22 2 11 15 2 nenh l=2e-07 w=1.1e-06 
+ as=5.76399e-13 ad=1.30942e-12 ps=1.98e-06 pd=4.01923e-06 
+ nrs=0.476363 nrd=1.08216 
md23 2 4 3 2 nenh l=2e-07 w=1.1e-06 
+ as=4.58333e-13 ad=1.30942e-12 ps=1.34444e-06 pd=4.01923e-06 
+ nrs=0.378788 nrd=1.08216 
c40 2 9 3.0125e-13
c41 2 3 5.6252e-14
c42 2 7 1.9336e-13
c43 2 8 3.68023e-13
c44 2 15 1.43756e-13
c45 2 5 1.9336e-13
c46 2 6 2.86102e-13
c47 14 2 3.7502e-14
c48 1 2 8.7375e-14
c49 2 13 2.38125e-13
c50 2 4 1.60877e-13
c51 2 12 2.38125e-13
c52 2 11 1.42127e-13
c53 15 10 5.3125e-14
c54 5 10 2.1e-14
c55 12 11 1.6632e-14
c56 6 10 2.9e-14
c57 11 15 2.1255e-14
c58 11 5 2.8508e-14
c59 7 13 3.1632e-14
c60 12 15 1.188e-14
c61 12 5 3.1632e-14
c62 4 7 2.8508e-14
c63 12 6 2.4948e-14
c64 13 9 4.752e-15
c65 15 5 9.1125e-14
c66 8 13 2.4948e-14
c67 4 9 6.627e-15
c68 7 10 2.1e-14
c69 3 7 9.1125e-14
c70 9 10 5.625e-14
c71 8 10 2.1e-14
c72 3 9 1.875e-15
c73 14 6 6e-14
c74 11 9 6.627e-15
c75 12 9 4.752e-15
c76 15 9 1.875e-15
c77 5 9 1.5e-14
c78 15 8 8.38199e-14
c79 6 9 1.5e-14
c80 4 13 1.6632e-14
c81 7 9 1.5e-14
c82 3 13 1.188e-14
c83 3 4 2.1255e-14
c84 8 9 1.5e-14
c85 1 6 3.8133e-14
c86 3 10 5.3125e-14
.ends FlashLatch
.subckt z2xFlashLatch 1 2 3 4 5
+ 6 7 8 9 10 11
+ 12 13 14
xFlashLatch#1 14 1 10 9 5
+ 6 3 4 12 2 FlashLatch
xFlashLatch#0 13 1 7 8 5
+ 6 3 4 11 2 FlashLatch
.ends z2xFlashLatch
.subckt z65xFlashLatch 1 2 3 4 5
+ 6 7 8 9 10 11
+ 12 13 14 15 16 17
+ 18 19 20 21 22 23
+ 24 25 26 27 28 29
+ 30 31 32 33 34 35
+ 36 37 38 39 40 41
+ 42 43 44 45 46 47
+ 48 49 50 51 52 53
+ 54 55 56 57 58 59
+ 60 61 62 63 64 65
+ 66 67 68 69 70 71
+ 72 73 74 75 76 77
+ 78 79 80 81 82 83
+ 84 85 86 87 88 89
+ 90 91 92 93 94 95
+ 96 97 98 99 100 101
+ 102 103 104 105 106 107
+ 108 109 110 111 112 113
+ 114 115 116 117 118 119
+ 120 121 122 123 124 125
+ 126 127 128 129 130 131
+ 132 133 134 135 136 137
+ 138 139 140 141 142 143
+ 144 145 146 147 148 149
+ 150 151 152 153 154 155
+ 156 157 158 159 160 161
+ 162 163 164 165 166 167
+ 168 169 170 171 172 173
+ 174 175 176 177 178 179
+ 180 181 182 183 184 185
+ 186 187 188 189 190 191
+ 192 193 194 195 196 197
+ 198 199 200 201 202 203
+ 204 205 206 207 208 209
+ 210 211 212 213 214 215
+ 216 217 218 219 220 221
+ 222 223 224 225 226 227
+ 228 229 230 231 232 233
+ 234 235 236 237 238 239
+ 240 241 242 243 244 245
+ 246 247 248 249 250 251
+ 252 253 254 255 256 257
+ 258 259 260 261 262 263
+ 264 265 266
xFlashLatch#0 195 1 101 87 145
+ 156 123 134 142 2 FlashLatch
xz2xFlashLatch#0#0 1 2 123 134 145
+ 156 33 266 216 34 256
+ 225 129 192 z2xFlashLatch
xz2xFlashLatch#0#1 1 2 123 134 145
+ 156 27 260 203 239 221
+ 238 160 140 z2xFlashLatch
xz2xFlashLatch#0#2 1 2 123 134 145
+ 156 71 54 16 38 98
+ 75 183 141 z2xFlashLatch
xz2xFlashLatch#0#3 1 2 123 134 145
+ 156 106 92 65 79 21
+ 237 191 170 z2xFlashLatch
xz2xFlashLatch#0#4 1 2 123 134 145
+ 156 232 197 200 233 122
+ 113 137 188 z2xFlashLatch
xz2xFlashLatch#0#5 1 2 123 134 145
+ 156 223 7 13 36 74
+ 47 139 194 z2xFlashLatch
xz2xFlashLatch#0#6 1 2 123 134 145
+ 156 31 264 213 248 236
+ 11 169 152 z2xFlashLatch
xz2xFlashLatch#0#7 1 2 123 134 145
+ 156 73 58 22 42 112
+ 93 187 153 z2xFlashLatch
xz2xFlashLatch#0#8 1 2 123 134 145
+ 156 107 95 69 83 48
+ 10 193 180 z2xFlashLatch
xz2xFlashLatch#0#9 1 2 123 134 145
+ 156 242 205 209 245 212
+ 227 150 190 z2xFlashLatch
xz2xFlashLatch#0#10 1 2 123 134 145
+ 156 229 167 109 117 105
+ 108 146 173 z2xFlashLatch
xz2xFlashLatch#0#11 1 2 123 134 145
+ 156 28 261 204 240 86
+ 199 174 128 z2xFlashLatch
xz2xFlashLatch#0#12 1 2 123 134 145
+ 156 263 234 243 3 259
+ 210 144 159 z2xFlashLatch
xz2xFlashLatch#0#13 1 2 123 134 145
+ 156 57 37 39 60 8
+ 26 172 125 z2xFlashLatch
xz2xFlashLatch#0#14 1 2 123 134 145
+ 156 94 78 80 96 62
+ 30 126 155 z2xFlashLatch
xz2xFlashLatch#0#15 1 2 123 134 145
+ 156 224 110 111 118 207
+ 77 157 182 z2xFlashLatch
xz2xFlashLatch#0#16 1 2 123 134 145
+ 156 32 265 214 198 226
+ 249 124 138 z2xFlashLatch
xz2xFlashLatch#0#17 1 2 123 134 145
+ 156 5 246 250 9 29
+ 253 154 168 z2xFlashLatch
xz2xFlashLatch#0#18 1 2 123 134 145
+ 156 61 41 43 63 40
+ 53 181 135 z2xFlashLatch
xz2xFlashLatch#0#19 1 2 123 134 145
+ 156 97 82 84 99 81
+ 55 136 165 z2xFlashLatch
xz2xFlashLatch#0#20 1 2 123 134 145
+ 156 230 178 114 119 252
+ 196 166 186 z2xFlashLatch
xz2xFlashLatch#0#21 1 2 123 134 145
+ 156 201 6 219 206 262
+ 18 133 151 z2xFlashLatch
xz2xFlashLatch#0#22 1 2 123 134 145
+ 156 14 251 254 17 56
+ 25 164 179 z2xFlashLatch
xz2xFlashLatch#0#23 1 2 123 134 145
+ 156 64 45 46 66 189
+ 72 185 148 z2xFlashLatch
xz2xFlashLatch#0#24 1 2 123 134 145
+ 156 100 85 88 102 218
+ 231 149 176 z2xFlashLatch
xz2xFlashLatch#0#25 1 2 123 134 145
+ 156 235 202 115 120 24
+ 244 177 132 z2xFlashLatch
xz2xFlashLatch#0#26 1 2 123 134 145
+ 156 208 15 222 215 35
+ 44 147 163 z2xFlashLatch
xz2xFlashLatch#0#27 1 2 123 134 145
+ 156 19 255 258 23 76
+ 51 175 130 z2xFlashLatch
xz2xFlashLatch#0#28 1 2 123 134 145
+ 156 67 49 52 70 241
+ 91 131 161 z2xFlashLatch
xz2xFlashLatch#0#29 1 2 123 134 145
+ 156 103 89 90 104 257
+ 4 162 184 z2xFlashLatch
xz2xFlashLatch#0#30 1 2 123 134 145
+ 156 247 211 116 121 50
+ 12 127 143 z2xFlashLatch
xz2xFlashLatch#0#31 1 2 123 134 145
+ 156 217 20 228 220 59
+ 68 158 171 z2xFlashLatch
.ends z65xFlashLatch
.subckt FlashOFlo 1 2 3 4 5
md24 6 4 2 2 nenh l=2e-07 w=3.1e-06 
+ as=3.04745e-12 ad=7.8288e-13 ps=6.88304e-06 pd=6.8305e-07 
+ nrs=0.317113 nrd=0.0814651 
md25 2 7 3 2 nenh l=2e-07 w=1.4e-06 
+ as=6.29999e-13 ad=1.37627e-12 ps=9e-07 pd=3.10847e-06 
+ nrs=0.321428 nrd=0.702178 
md26 3 7 2 2 nenh l=2e-07 w=1.4e-06 
+ as=1.37627e-12 ad=6.29999e-13 ps=3.10847e-06 pd=9e-07 
+ nrs=0.702178 nrd=0.321428 
md27 7 1 6 2 nenh l=2e-07 w=2.8e-06 
+ as=7.07117e-13 ad=1.54e-12 ps=6.16948e-07 pd=4.39999e-06 
+ nrs=0.0901935 nrd=0.196429 
md28 7 4 5 5 penh l=2e-07 w=1.5e-06 
+ as=1.85281e-12 ad=7.99999e-13 ps=4.07745e-06 pd=3.1e-06 
+ nrs=0.823473 nrd=0.355556 
md29 5 7 3 5 penh l=2e-07 w=2.8e-06 
+ as=1.26e-12 ad=3.45858e-12 ps=9e-07 pd=7.61127e-06 
+ nrs=0.160714 nrd=0.441146 
md30 3 7 5 5 penh l=2e-07 w=2.8e-06 
+ as=3.45858e-12 ad=1.26e-12 ps=7.61127e-06 pd=9e-07 
+ nrs=0.441146 nrd=0.160714 
c87 2 3 3.89625e-13
c88 2 7 5.20127e-13
c89 1 2 1.74e-13
c90 2 4 3.51567e-13
c91 7 5 2.36877e-13
c92 6 5 5.5875e-14
c93 3 5 5.625e-15
c94 1 5 9.8823e-14
c95 2 5 4.90625e-13
c96 4 5 5.675e-14
c97 3 7 4.6332e-14
c98 1 7 1.4256e-14
.ends FlashOFlo
.subckt Flash3ANDS 1 2 3 4 5
+ 6 7 8 9
md31 9 3 10 9 penh l=1.1e-06 w=5e-07 
+ as=3.47499e-13 ad=4.78289e-13 ps=1.45e-06 pd=1.26316e-06 
+ nrs=1.39 nrd=1.91316 
md32 10 7 9 9 penh l=2e-07 w=1.5e-06 
+ as=1.43487e-12 ad=1.0425e-12 ps=3.78947e-06 pd=4.35e-06 
+ nrs=0.637719 nrd=0.463333 
md33 9 10 3 9 penh l=2e-07 w=2.8e-06 
+ as=1.26e-12 ad=2.67841e-12 ps=9e-07 pd=7.07368e-06 
+ nrs=0.160714 nrd=0.341635 
md34 3 10 9 9 penh l=2e-07 w=2.8e-06 
+ as=2.67841e-12 ad=1.26e-12 ps=7.07368e-06 pd=9e-07 
+ nrs=0.341635 nrd=0.160714 
md35 10 2 11 4 nenh l=2e-07 w=2.8e-06 
+ as=6.99999e-13 ad=1.54e-12 ps=5e-07 pd=4.39999e-06 
+ nrs=0.0892856 nrd=0.196429 
md36 12 7 4 4 nenh l=2e-07 w=3.1e-06 
+ as=2.79e-12 ad=7.8288e-13 ps=6.14745e-06 pd=6.8305e-07 
+ nrs=0.290322 nrd=0.0814651 
md37 4 10 3 4 nenh l=2e-07 w=1.4e-06 
+ as=6.29999e-13 ad=1.26e-12 ps=9e-07 pd=2.77627e-06 
+ nrs=0.321428 nrd=0.642857 
md38 3 10 4 4 nenh l=2e-07 w=1.4e-06 
+ as=1.26e-12 ad=6.29999e-13 ps=2.77627e-06 pd=9e-07 
+ nrs=0.642857 nrd=0.321428 
md39 13 1 12 4 nenh l=2e-07 w=2.8e-06 
+ as=7.07117e-13 ad=6.99999e-13 ps=6.16948e-07 pd=5e-07 
+ nrs=0.0901935 nrd=0.0892856 
md40 11 5 13 4 nenh l=2e-07 w=2.8e-06 
+ as=6.99999e-13 ad=6.99999e-13 ps=5e-07 pd=5e-07 
+ nrs=0.0892856 nrd=0.0892856 
c99 4 8 2.8875e-13
c100 2 4 1.3034e-13
c101 4 5 2.6558e-13
c102 3 4 5.79e-13
c103 4 6 2.66375e-13
c104 1 4 1.16e-13
c105 10 4 5.29754e-13
c106 4 7 3.15307e-13
c107 7 9 5.075e-14
c108 11 6 1.25e-14
c109 3 10 7.722e-14
c110 11 9 4.5e-14
c111 12 6 1.4375e-14
c112 3 9 3.75e-15
c113 5 6 1.188e-14
c114 1 5 1.188e-14
c115 6 8 1.782e-14
c116 1 8 1.782e-14
c117 12 9 4.725e-14
c118 10 8 3.126e-14
c119 5 9 1.07375e-13
c120 5 7 5.8076e-14
c121 13 6 1.25e-14
c122 8 9 1.68125e-13
c123 7 8 2.688e-14
c124 1 6 1.188e-14
c125 13 9 4.5e-14
c126 10 6 4.314e-14
c127 1 10 1.5444e-14
c128 2 6 1.188e-14
c129 3 8 2.8125e-14
c130 6 9 1.61698e-13
c131 1 9 7.5012e-14
c132 6 7 4.47e-14
c133 4 9 3.9725e-13
c134 10 9 1.75377e-13
c135 2 9 2.1e-14
.ends Flash3ANDS
.subckt z2xFlashANDN 1 2 3 4 5
+ 6 7 8 9
xFlashOFlo#0 4 1 8 7 2 FlashOFlo
xFlash3ANDS#0 2 3 9 1 5
+ 4 7 6 2 Flash3ANDS
.ends z2xFlashANDN
.subckt Flash3ANDN 1 2 3 4 5
+ 6 7 8 9
md41 10 7 4 4 nenh l=2e-07 w=3.1e-06 
+ as=2.79e-12 ad=7.8288e-13 ps=6.14745e-06 pd=6.8305e-07 
+ nrs=0.290322 nrd=0.0814651 
md42 4 11 3 4 nenh l=2e-07 w=1.4e-06 
+ as=6.29999e-13 ad=1.26e-12 ps=9e-07 pd=2.77627e-06 
+ nrs=0.321428 nrd=0.642857 
md43 3 11 4 4 nenh l=2e-07 w=1.4e-06 
+ as=1.26e-12 ad=6.29999e-13 ps=2.77627e-06 pd=9e-07 
+ nrs=0.642857 nrd=0.321428 
md44 12 1 10 4 nenh l=2e-07 w=2.8e-06 
+ as=7.07117e-13 ad=6.99999e-13 ps=6.16948e-07 pd=5e-07 
+ nrs=0.0901935 nrd=0.0892856 
md45 13 5 12 4 nenh l=2e-07 w=2.8e-06 
+ as=6.99999e-13 ad=6.99999e-13 ps=5e-07 pd=5e-07 
+ nrs=0.0892856 nrd=0.0892856 
md46 11 2 13 4 nenh l=2e-07 w=2.8e-06 
+ as=6.99999e-13 ad=1.54e-12 ps=5e-07 pd=4.39999e-06 
+ nrs=0.0892856 nrd=0.196429 
md47 9 3 11 9 penh l=1.1e-06 w=5e-07 
+ as=4.09999e-13 ad=5.7763e-13 ps=1.7e-06 pd=1.27631e-06 
+ nrs=1.64 nrd=2.31052 
md48 11 7 9 9 penh l=2e-07 w=1.5e-06 
+ as=1.73289e-12 ad=1.23e-12 ps=3.82894e-06 pd=5.1e-06 
+ nrs=0.770174 nrd=0.546666 
md49 9 11 3 9 penh l=2e-07 w=2.8e-06 
+ as=1.26e-12 ad=3.23473e-12 ps=9e-07 pd=7.14736e-06 
+ nrs=0.160714 nrd=0.412594 
md50 3 11 9 9 penh l=2e-07 w=2.8e-06 
+ as=3.23473e-12 ad=1.26e-12 ps=7.14736e-06 pd=9e-07 
+ nrs=0.412594 nrd=0.160714 
c136 4 8 2.56875e-13
c137 3 4 5.38e-13
c138 11 4 5.33629e-13
c139 2 4 1.28e-13
c140 4 5 2.74375e-13
c141 4 7 3.16623e-13
c142 4 6 3.3484e-13
c143 1 4 8.658e-14
c144 6 9 9.3e-14
c145 2 8 1.782e-14
c146 5 8 1.782e-14
c147 7 9 5.075e-14
c148 11 8 3.56349e-14
c149 6 7 4.47e-14
c150 13 9 4.5e-14
c151 13 6 1.25e-14
c152 3 8 6.7329e-14
c153 1 9 2.1e-14
c154 1 6 1.188e-14
c155 2 11 1.782e-14
c156 11 5 1.782e-14
c157 8 9 1.75e-13
c158 7 8 2.688e-14
c159 3 11 6.2964e-14
c160 10 9 4.725e-14
c161 2 9 7.1073e-14
c162 10 6 1.4375e-14
c163 2 6 1.188e-14
c164 5 9 1.45012e-13
c165 5 6 1.188e-14
c166 11 9 2.19127e-13
c167 4 9 4.26125e-13
c168 11 6 2.532e-14
c169 5 7 5.8076e-14
c170 3 9 4.0625e-14
c171 12 9 4.5e-14
c172 12 6 1.25e-14
.ends Flash3ANDN
.subckt z2xFlash3AND 1 2 3 4 5
+ 6 7 8 9 10 11
+ 12 13
xFlash3ANDN#0 6 4 13 1 5
+ 9 7 10 2 Flash3ANDN
xFlash3ANDS#0 5 8 11 1 3
+ 4 7 12 2 Flash3ANDS
.ends z2xFlash3AND
.subckt FlashUFlo 1 2 3 4 5
+ 6 7 8
md51 8 7 9 8 penh l=1.1e-06 w=5e-07 
+ as=3.47499e-13 ad=4.78289e-13 ps=1.45e-06 pd=1.26316e-06 
+ nrs=1.39 nrd=1.91316 
md52 9 5 8 8 penh l=2e-07 w=1.5e-06 
+ as=1.43487e-12 ad=1.0425e-12 ps=3.78947e-06 pd=4.35e-06 
+ nrs=0.637719 nrd=0.463333 
md53 8 9 7 8 penh l=2e-07 w=2.8e-06 
+ as=1.26e-12 ad=2.67841e-12 ps=9e-07 pd=7.07368e-06 
+ nrs=0.160714 nrd=0.341635 
md54 7 9 8 8 penh l=2e-07 w=2.8e-06 
+ as=2.67841e-12 ad=1.26e-12 ps=7.07368e-06 pd=9e-07 
+ nrs=0.341635 nrd=0.160714 
md55 9 3 10 2 nenh l=2e-07 w=2.8e-06 
+ as=6.99999e-13 ad=1.54e-12 ps=5e-07 pd=4.39999e-06 
+ nrs=0.0892856 nrd=0.196429 
md56 11 5 2 2 nenh l=2e-07 w=3.1e-06 
+ as=3.04745e-12 ad=7.8288e-13 ps=6.88304e-06 pd=6.8305e-07 
+ nrs=0.317113 nrd=0.0814651 
md57 2 9 7 2 nenh l=2e-07 w=1.4e-06 
+ as=6.29999e-13 ad=1.37627e-12 ps=9e-07 pd=3.10847e-06 
+ nrs=0.321428 nrd=0.702178 
md58 7 9 2 2 nenh l=2e-07 w=1.4e-06 
+ as=1.37627e-12 ad=6.29999e-13 ps=3.10847e-06 pd=9e-07 
+ nrs=0.702178 nrd=0.321428 
md59 10 1 11 2 nenh l=2e-07 w=2.8e-06 
+ as=7.07117e-13 ad=6.99999e-13 ps=6.16948e-07 pd=5e-07 
+ nrs=0.0901935 nrd=0.0892856 
c173 2 6 2.8875e-13
c174 2 3 1.83e-13
c175 2 7 5.79e-13
c176 2 4 2.85125e-13
c177 1 2 1.16e-13
c178 2 9 5.51629e-13
c179 2 5 3.16623e-13
c180 5 6 2.688e-14
c181 11 4 1.4375e-14
c182 3 4 1.188e-14
c183 4 5 4.47e-14
c184 1 6 1.782e-14
c185 10 4 1.25e-14
c186 7 9 7.722e-14
c187 4 6 1.782e-14
c188 1 4 1.188e-14
c189 7 8 3.75e-15
c190 11 8 4.725e-14
c191 3 8 1.05125e-13
c192 2 8 3.9725e-13
c193 5 8 5.075e-14
c194 6 9 3.126e-14
c195 1 9 1.5444e-14
c196 10 8 4.5e-14
c197 6 8 1.68125e-13
c198 4 9 4.314e-14
c199 1 8 7.5012e-14
c200 4 8 1.61698e-13
c201 3 5 5.8076e-14
c202 6 7 2.8125e-14
c203 9 8 1.92877e-13
c204 1 3 1.188e-14
.ends FlashUFlo
.subckt z2xFlashANDS 1 2 3 4 5
+ 6 7 8 9 10 11
+ 12
xFlash3ANDN#0 5 4 11 1 8
+ 3 6 9 2 Flash3ANDN
xFlashUFlo#0 8 1 7 4 6
+ 10 12 2 FlashUFlo
.ends z2xFlashANDS
.subckt FlashOneHot 1 2 3 4 5
+ 6 7 8 9 10 11
+ 12 13 14 15 16 17
+ 18 19 20 21 22 23
+ 24 25 26 27 28 29
+ 30 31 32 33 34 35
+ 36 37 38 39 40 41
+ 42 43 44 45 46 47
+ 48 49 50 51 52 53
+ 54 55 56 57 58 59
+ 60 61 62 63 64 65
+ 66 67 68 69 70 71
+ 72 73 74 75 76 77
+ 78 79 80 81 82 83
+ 84 85 86 87 88 89
+ 90 91 92 93 94 95
+ 96 97 98 99 100 101
+ 102 103 104 105 106 107
+ 108 109 110 111 112 113
+ 114 115 116 117 118 119
+ 120 121 122 123 124 125
+ 126 127 128 129 130 131
+ 132 133 134 135 136 137
+ 138 139 140 141 142 143
+ 144 145 146 147 148 149
+ 150 151 152 153 154 155
+ 156 157 158 159 160 161
+ 162 163 164 165 166 167
+ 168 169 170 171 172 173
+ 174 175 176 177 178 179
+ 180 181 182 183 184 185
+ 186 187 188 189 190 191
+ 192 193 194 195 196 197
+ 198 199 200 201 202
xz65xFlashLatch#0 1 2 203 28 204
+ 205 206 29 207 30 31
+ 32 208 209 210 211 212
+ 33 213 214 34 215 216
+ 35 36 37 217 218 38
+ 39 219 220 221 222 40
+ 223 224 225 226 41 227
+ 228 229 42 230 231 43
+ 44 232 46 47 233 48
+ 234 49 50 235 236 51
+ 237 238 52 239 240 241
+ 242 243 53 244 245 246
+ 54 247 55 56 57 58
+ 248 249 250 59 251 252
+ 253 254 60 255 256 257
+ 258 61 259 62 260 261
+ 262 263 63 264 265 266
+ 267 268 269 64 270 271
+ 65 272 273 274 66 67
+ 275 276 277 278 279 280
+ 281 282 68 132 69 72
+ 74 75 77 78 80 83
+ 86 88 154 91 92 94
+ 95 96 97 99 45 100
+ 102 26 105 108 111 113
+ 115 118 119 121 124 125
+ 90 126 127 129 130 131
+ 134 136 141 143 144 283
+ 147 148 150 152 153 156
+ 157 158 160 161 284 163
+ 164 166 168 170 172 177
+ 179 180 181 3 192 193
+ 194 196 198 202 4 285
+ 286 5 287 288 289 290
+ 291 292 293 6 294 295
+ 7 296 8 297 298 299
+ 300 301 9 302 303 10
+ 304 305 306 11 12 13
+ 307 308 309 14 310 311
+ 312 313 15 16 17 314
+ 315 18 316 317 19 318
+ 319 320 321 20 322 323
+ 21 22 324 325 23 24
+ 326 25 327 328 27 329
+ 330 331 332 z65xFlashLatch
xz2xFlashANDN#0 1 2 307 255 266
+ 45 26 162 176 z2xFlashANDN
xz2xFlash3AND#0#0 1 2 217 327 314
+ 246 26 300 290 17 185
+ 10 137 z2xFlash3AND
xz2xFlash3AND#0#1 1 2 246 234 225
+ 270 26 290 211 56 106
+ 63 93 z2xFlash3AND
xz2xFlash3AND#0#2 1 2 270 259 249
+ 310 26 211 241 16 149
+ 34 73 z2xFlash3AND
xz2xFlash3AND#0#3 1 2 310 285 311
+ 305 26 241 287 67 103
+ 68 187 z2xFlash3AND
xz2xFlash3AND#0#4 1 2 305 206 223
+ 219 26 287 208 43 200
+ 55 138 z2xFlash3AND
xz2xFlash3AND#0#5 1 2 219 330 321
+ 247 26 208 297 31 184
+ 15 159 z2xFlash3AND
xz2xFlash3AND#0#6 1 2 247 236 228
+ 271 26 297 215 62 104
+ 66 122 z2xFlash3AND
xz2xFlash3AND#0#7 1 2 271 261 252
+ 316 26 215 244 30 167
+ 44 70 z2xFlash3AND
xz2xFlash3AND#0#8 1 2 316 292 318
+ 308 26 244 295 13 133
+ 8 186 z2xFlash3AND
xz2xFlash3AND#0#9 1 2 308 283 278
+ 218 26 295 272 65 87
+ 64 107 z2xFlash3AND
xz2xFlash3AND#0#10 1 2 218 328 315
+ 329 26 272 291 5 120
+ 60 195 z2xFlash3AND
xz2xFlash3AND#0#11 1 2 329 312 203
+ 235 26 291 317 7 71
+ 25 142 z2xFlash3AND
xz2xFlash3AND#0#12 1 2 235 224 237
+ 260 26 317 226 37 188
+ 29 165 z2xFlash3AND
xz2xFlash3AND#0#13 1 2 260 248 262
+ 306 26 226 250 39 110
+ 52 128 z2xFlash3AND
xz2xFlash3AND#0#14 1 2 306 273 279
+ 220 26 250 274 58 174
+ 6 76 z2xFlash3AND
xz2xFlash3AND#0#15 1 2 220 331 286
+ 204 26 274 298 20 139
+ 12 189 z2xFlash3AND
xz2xFlash3AND#0#16 1 2 204 319 207
+ 238 26 298 322 22 98
+ 38 112 z2xFlash3AND
xz2xFlash3AND#0#17 1 2 238 227 239
+ 263 26 322 229 48 169
+ 41 178 z2xFlash3AND
xz2xFlash3AND#0#18 1 2 263 251 264
+ 309 26 229 253 49 79
+ 59 145 z2xFlash3AND
xz2xFlash3AND#0#19 1 2 309 284 280
+ 288 26 253 275 4 183
+ 21 109 z2xFlash3AND
xz2xFlash3AND#0#20 1 2 288 205 293
+ 209 26 275 302 33 114
+ 27 171 z2xFlash3AND
xz2xFlash3AND#0#21 1 2 209 323 212
+ 240 26 302 324 36 123
+ 50 82 z2xFlash3AND
xz2xFlash3AND#0#22 1 2 240 230 242
+ 265 26 324 231 54 81
+ 3 191 z2xFlash3AND
xz2xFlash3AND#0#23 1 2 265 254 267
+ 313 26 231 256 14 199
+ 9 116 z2xFlash3AND
xz2xFlash3AND#0#24 1 2 313 289 281
+ 294 26 256 276 19 173
+ 35 135 z2xFlash3AND
xz2xFlash3AND#0#25 1 2 294 210 299
+ 213 26 276 304 42 84
+ 40 89 z2xFlash3AND
xz2xFlash3AND#0#26 1 2 213 325 216
+ 243 26 304 326 47 146
+ 57 201 z2xFlash3AND
xz2xFlash3AND#0#27 1 2 243 232 245
+ 268 26 326 233 61 101
+ 18 175 z2xFlash3AND
xz2xFlash3AND#0#28 1 2 268 257 269
+ 320 26 233 258 28 197
+ 24 85 z2xFlash3AND
xz2xFlash3AND#0#29 1 2 320 296 282
+ 301 26 258 277 32 151
+ 46 155 z2xFlash3AND
xz2xFlash3AND#0#30 1 2 301 214 303
+ 266 26 277 307 53 190
+ 51 117 z2xFlash3AND
xz2xFlashANDS#0 1 2 300 332 217
+ 26 221 222 11 23 140
+ 182
+ z2xFlashANDS
.ends FlashOneHot
.subckt ConvertLatch 1 2 3 4 5
+ 6 7 8
md60 8 4 2 8 penh l=2e-07 w=2.1e-06 
+ as=9.44999e-13 ad=2.00973e-12 ps=9e-07 pd=4.6421e-06 
+ nrs=0.214286 nrd=0.455722 
md61 2 4 8 8 penh l=2e-07 w=2.1e-06 
+ as=2.00973e-12 ad=9.44999e-13 ps=4.6421e-06 pd=9e-07 
+ nrs=0.455722 nrd=0.214286 
md62 9 2 8 8 penh l=2e-07 w=1.4e-06 
+ as=1.33982e-12 ad=5.59999e-13 ps=3.09473e-06 pd=1.66666e-06 
+ nrs=0.683583 nrd=0.285714 
md63 10 11 8 8 penh l=2e-07 w=2.7e-06 
+ as=2.77534e-12 ad=9.87803e-13 ps=6.41052e-06 pd=1.28049e-06 
+ nrs=0.330005 nrd=0.158049 
md64 1 12 8 8 penh l=2e-07 w=2.7e-06 
+ as=2.77534e-12 ad=1.01e-12 ps=6.41052e-06 pd=2.9e-06 
+ nrs=0.330005 nrd=0.1616 
md65 11 4 9 3 nenh l=2e-07 w=7e-07 
+ as=3.15e-13 ad=5.59999e-13 ps=9e-07 pd=2.3e-06 
+ nrs=0.642857 nrd=1.14286 
md66 9 2 3 3 nenh l=2e-07 w=7e-07 
+ as=1.498e-12 ad=3.15e-13 ps=3.18e-06 pd=9e-07 
+ nrs=3.05714 nrd=0.642857 
md67 11 5 9 8 penh l=2e-07 w=7e-07 
+ as=2.8e-13 ad=5.59999e-13 ps=8.33332e-07 pd=2.3e-06 
+ nrs=0.571428 nrd=1.14286 
md68 10 11 3 3 nenh l=2e-07 w=1.4e-06 
+ as=2.99599e-12 ad=6.29999e-13 ps=6.35999e-06 pd=9e-07 
+ nrs=1.52857 nrd=0.321428 
md69 1 12 3 3 nenh l=2e-07 w=1.4e-06 
+ as=2.99599e-12 ad=1.12e-12 ps=6.35999e-06 pd=3e-06 
+ nrs=1.52857 nrd=0.571428 
md70 12 6 10 3 nenh l=2e-07 w=1.4e-06 
+ as=6.29999e-13 ad=1.12e-12 ps=9e-07 pd=3e-06 
+ nrs=0.321428 nrd=0.571428 
md71 10 7 12 8 penh l=2e-07 w=1.6e-06 
+ as=8.29999e-13 ad=6.32194e-13 ps=3.2e-06 pd=8.19511e-07 
+ nrs=0.324219 nrd=0.246951 
c205 3 4 5.39025e-13
c206 1 3 4.18752e-13
c207 12 3 1.6275e-13
c208 10 3 6.2502e-14
c209 3 6 1.54199e-13
c210 3 7 3.48318e-13
c211 11 3 3.57875e-13
c212 3 5 1.58431e-13
c213 9 3 4.375e-14
c214 2 3 9.54e-13
c215 2 4 5.8512e-14
c216 12 10 2.0625e-14
c217 12 7 9.504e-15
c218 12 8 2.875e-14
c219 6 7 4.5e-15
c220 5 8 3.75e-14
c221 12 11 4.752e-15
c222 1 8 1.4725e-13
c223 10 7 1.188e-14
c224 12 2 1.188e-14
c225 6 8 2.1e-14
c226 2 5 3.75e-15
c227 11 6 6.75e-15
c228 1 2 3.75e-14
c229 2 6 1.5e-14
c230 9 5 4.5e-15
c231 7 8 8.7528e-14
c232 1 4 3.87599e-14
c233 11 7 6.75e-15
c234 2 7 1.5e-14
c235 4 8 1.57877e-13
c236 2 8 1.20625e-13
c237 11 4 1.5e-14
c238 3 8 3.06e-13
c239 11 2 5.7024e-14
c240 12 1 1.188e-14
.ends ConvertLatch
.subckt z2xConvertLatch 1 2 3 4 5
+ 6 7 8 9 10
xConvertLatch#0 4 7 1 5 3
+ 6 9 2 ConvertLatch
xConvertLatch#1 8 10 1 5 3
+ 6 9 2 ConvertLatch
.ends z2xConvertLatch
.subckt z7xConvertLatch 1 2 3 4 5
+ 6 7 8 9 10 11
+ 12 13 14 15 16 17
+ 18 19 20
xz2xConvertLatch#0#0 1 2 4 7 3
+ 5 9 16 6 12 z2xConvertLatch
xz2xConvertLatch#0#1 1 2 4 10 3
+ 5 15 17 6 18 z2xConvertLatch
xz2xConvertLatch#0#2 1 2 4 11 3
+ 5 14 8 6 19 z2xConvertLatch
xConvertLatch#0 13 20 1 3 4
+ 5 6 2 ConvertLatch
.ends z7xConvertLatch
.subckt AtoDRtgW 1 2 3 4 5
c241 1 4 8.37177e-11
c242 2 4 2.99996e-12
c243 3 4 2.71743e-12
c244 1 3 1.92e-12
c245 1 2 2.4e-13
c246 2 3 3.2e-14
.ends AtoDRtgW
.subckt CDLabels 1 2 3 4 5
+ 6 7 8 9 10 11
+ 12 13 14 15 16 17
+ 18 19 20 21 22 23
+ 24 25 26 27 28 29
+ 30 31 32 33 34 35
+ 36 37 38 39 40 41
+ 42 43 44 45 46 47
+ 48 49 50 51 52 53
+ 54 55 56 57 58 59
+ 60 61 62 63 64 65
+ 66 67 68 69 70 71
+ 72 73 74 75 76 77
+ 78 79 80 81 82 83
+ 84 85 86 87 88 89
+ 90 91 92 93 94 95
+ 96 97 98 99 100 101
+ 102 103 104 105 106 107
+ 108 109 110 111 112 113
+ 114 115 116 117 118 119
+ 120 121 122 123 124 125
+ 126 127 128 129 130 131
+ 132 133 134 135 136 137
+ 138 139 140 141 142 143
+ 144 145 146 147 148 149
+ 150 151 152 153 154 155
+ 156 157 158 159 160 161
+ 162 163 164 165 166 167
c247 1 99 3.0625e-14
c248 99 166 3.0625e-14
c249 99 101 2.1875e-14
c250 99 103 2.1875e-14
c251 35 99 3.0625e-14
c252 9 99 3.0625e-14
c253 46 99 3.0625e-14
c254 99 114 2.1875e-14
c255 99 125 2.1875e-14
c256 57 99 3.0625e-14
c257 20 99 3.0625e-14
c258 68 99 3.0625e-14
c259 99 136 2.1875e-14
c260 99 147 2.1875e-14
c261 79 99 3.0625e-14
c262 31 99 3.0625e-14
c263 90 99 3.0625e-14
c264 99 158 2.1875e-14
c265 99 162 2.1875e-14
c266 95 99 3.0625e-14
c267 3 99 3.0625e-14
c268 96 99 3.0625e-14
c269 99 163 2.1875e-14
c270 99 164 2.1875e-14
c271 97 99 3.0625e-14
c272 4 99 3.0625e-14
c273 98 99 3.0625e-14
c274 99 165 2.1875e-14
c275 99 104 2.1875e-14
c276 36 99 3.0625e-14
c277 5 99 3.0625e-14
c278 37 99 3.0625e-14
c279 99 105 2.1875e-14
c280 99 106 2.1875e-14
c281 38 99 3.0625e-14
c282 6 99 3.0625e-14
c283 39 99 3.0625e-14
c284 99 107 2.1875e-14
c285 99 108 2.1875e-14
c286 40 99 3.0625e-14
c287 7 99 3.0625e-14
c288 41 99 3.0625e-14
c289 99 109 2.1875e-14
c290 99 110 2.1875e-14
c291 42 99 3.0625e-14
c292 8 99 3.0625e-14
c293 43 99 3.0625e-14
c294 99 111 2.1875e-14
c295 99 112 2.1875e-14
c296 44 99 3.0625e-14
c297 10 99 3.0625e-14
c298 45 99 3.0625e-14
c299 99 113 2.1875e-14
c300 99 115 2.1875e-14
c301 47 99 3.0625e-14
c302 11 99 3.0625e-14
c303 48 99 3.0625e-14
c304 99 116 2.1875e-14
c305 99 117 2.1875e-14
c306 49 99 3.0625e-14
c307 12 99 3.0625e-14
c308 50 99 3.0625e-14
c309 99 118 2.1875e-14
c310 99 119 2.1875e-14
c311 51 99 3.0625e-14
c312 13 99 3.0625e-14
c313 52 99 3.0625e-14
c314 99 120 2.1875e-14
c315 99 121 2.1875e-14
c316 53 99 3.0625e-14
c317 14 99 3.0625e-14
c318 54 99 3.0625e-14
c319 99 122 2.1875e-14
c320 99 123 2.1875e-14
c321 55 99 3.0625e-14
c322 15 99 3.0625e-14
c323 56 99 3.0625e-14
c324 99 124 2.1875e-14
c325 99 126 2.1875e-14
c326 58 99 3.0625e-14
c327 16 99 3.0625e-14
c328 59 99 3.0625e-14
c329 99 127 2.1875e-14
c330 99 128 2.1875e-14
c331 60 99 3.0625e-14
c332 17 99 3.0625e-14
c333 61 99 3.0625e-14
c334 99 129 2.1875e-14
c335 99 130 2.1875e-14
c336 62 99 3.0625e-14
c337 18 99 3.0625e-14
c338 63 99 3.0625e-14
c339 99 131 2.1875e-14
c340 99 132 2.1875e-14
c341 64 99 3.0625e-14
c342 19 99 3.0625e-14
c343 65 99 3.0625e-14
c344 99 133 2.1875e-14
c345 99 134 2.1875e-14
c346 66 99 3.0625e-14
c347 21 99 3.0625e-14
c348 67 99 3.0625e-14
c349 99 135 2.1875e-14
c350 99 137 2.1875e-14
c351 69 99 3.0625e-14
c352 22 99 3.0625e-14
c353 70 99 3.0625e-14
c354 99 138 2.1875e-14
c355 99 139 2.1875e-14
c356 71 99 3.0625e-14
c357 23 99 3.0625e-14
c358 72 99 3.0625e-14
c359 99 140 2.1875e-14
c360 99 141 2.1875e-14
c361 73 99 3.0625e-14
c362 24 99 3.0625e-14
c363 74 99 3.0625e-14
c364 99 142 2.1875e-14
c365 99 143 2.1875e-14
c366 75 99 3.0625e-14
c367 25 99 3.0625e-14
c368 76 99 3.0625e-14
c369 99 144 2.1875e-14
c370 99 145 2.1875e-14
c371 77 99 3.0625e-14
c372 26 99 3.0625e-14
c373 78 99 3.0625e-14
c374 99 146 2.1875e-14
c375 99 148 2.1875e-14
c376 80 99 3.0625e-14
c377 27 99 3.0625e-14
c378 81 99 3.0625e-14
c379 99 149 2.1875e-14
c380 99 150 2.1875e-14
c381 82 99 3.0625e-14
c382 28 99 3.0625e-14
c383 83 99 3.0625e-14
c384 99 151 2.1875e-14
c385 99 152 2.1875e-14
c386 84 99 3.0625e-14
c387 29 99 3.0625e-14
c388 85 99 3.0625e-14
c389 99 153 2.1875e-14
c390 99 154 2.1875e-14
c391 86 99 3.0625e-14
c392 30 99 3.0625e-14
c393 87 99 3.0625e-14
c394 99 155 2.1875e-14
c395 99 156 2.1875e-14
c396 88 99 3.0625e-14
c397 32 99 3.0625e-14
c398 89 99 3.0625e-14
c399 99 157 2.1875e-14
c400 99 159 2.1875e-14
c401 91 99 3.0625e-14
c402 33 99 3.0625e-14
c403 92 99 3.0625e-14
c404 99 160 2.1875e-14
c405 99 161 2.1875e-14
c406 93 99 3.0625e-14
c407 34 99 3.0625e-14
c408 94 99 3.0625e-14
c409 99 102 2.1875e-14
c410 99 100 3.0625e-14
c411 2 99 3.0625e-14
.ends CDLabels
.subckt ConvertDecode1 1 2 3 4 5
+ 6
md72 1 2 3 5 nenh l=2e-07 w=2.5e-06 
+ as=1.125e-12 ad=2e-12 ps=9e-07 pd=4.1e-06 
+ nrs=0.18 nrd=0.32 
md73 3 2 1 5 nenh l=2e-07 w=2.5e-06 
+ as=2e-12 ad=1.125e-12 ps=4.1e-06 pd=9e-07 
+ nrs=0.32 nrd=0.18 
c412 4 5 9.0625e-14
c413 3 5 1.66707e-13
c414 1 5 1.18125e-13
c415 2 5 1.99e-13
c416 2 3 2.975e-14
c417 1 3 2.45e-14
c418 3 4 1.75e-14
.ends ConvertDecode1
.subckt ConvertDecode0 1 2 3 4 5
+ 6
c419 4 5 1.33224e-13
c420 3 5 1.26875e-13
c421 2 5 9.0625e-14
c422 1 5 6.5625e-14
c423 1 4 2.45e-14
c424 3 4 2.45e-14
c425 2 4 1.75e-14
.ends ConvertDecode0
.subckt ConvertDecode 1 2 3 4 5
+ 6 7 8 9 10 11
+ 12 13 14 15 16 17
+ 18 19 20 21 22 23
+ 24 25 26 27 28 29
+ 30 31 32 33 34 35
+ 36 37 38 39 40 41
+ 42 43 44 45 46 47
+ 48 49 50 51 52 53
+ 54 55 56 57 58 59
+ 60 61 62 63 64 65
+ 66 67 68 69 70 71
+ 72 73 74 75 76 77
+ 78 79 80 81 82 83
+ 84 85 86 87 88 89
+ 90 91 92 93 94 95
+ 96 97 98 99 100 101
+ 102 103 104 105 106 107
+ 108 109 110 111 112 113
+ 114 115 116 117 118 119
+ 120 121 122 123 124 125
+ 126 127 128 129 130 131
+ 132 133 134 135 136 137
+ 138 139 140
xCDLables#0 1 1 1 1 1
+ 1 1 1 1 1 1
+ 1 1 1 1 1 1
+ 1 1 1 1 1 1
+ 1 1 1 1 1 1
+ 1 1 1 1 1 74
+ 72 115 86 42 57 94
+ 6 66 117 27 116 45
+ 56 131 7 76 120 91
+ 48 63 102 70 11 73
+ 121 35 49 96 109 12
+ 78 112 43 47 52 98
+ 61 15 14 123 137 53
+ 100 32 67 18 29 79
+ 140 38 103 132 20 83
+ 82 84 122 54 105 8
+ 41 118 138 1 89 37
+ 25 22 4 44 59 134
+ 34 88 95 9 24 108
+ 19 128 21 5 114 124
+ 46 65 129 3 68 31
+ 106 23 33 87 125 77
+ 60 107 133 17 99 80
+ 50 62 40 93 90 97
+ 16 28 126 130 30 71
+ 81 139 58 104 111 13
+ 55 119 10 135 39 92
+ 75 113 136 36 110 2 CDLabels
xDec#65#0 1 89 26 141 1
+ 2
+ ConvertDecode1
xDec#65#1 1 89 51 141 1
+ 2
+ ConvertDecode1
xDec#65#2 1 89 69 141 1
+ 2
+ ConvertDecode1
xDec#65#3 1 89 85 141 1
+ 2
+ ConvertDecode1
xDec#65#4 1 89 64 141 1
+ 2
+ ConvertDecode1
xDec#65#5 1 89 101 141 1
+ 2
+ ConvertDecode1
xDec#65#6 1 89 127 141 1
+ 2
+ ConvertDecode1
xDec#64#0 1 105 26 25 1
+ 2
+ ConvertDecode1
xDec#64#1 1 105 51 25 1
+ 2
+ ConvertDecode1
xDec#64#2 1 105 69 25 1
+ 2
+ ConvertDecode1
xDec#64#3 1 105 85 25 1
+ 2
+ ConvertDecode1
xDec#64#4 1 105 64 25 1
+ 2
+ ConvertDecode1
xDec#64#5 1 105 101 25 1
+ 2
+ ConvertDecode1
xDec#64#6 1 25 105 127 1
+ 2
+ ConvertDecode0
xDec#63#0 1 92 54 26 1
+ 2
+ ConvertDecode0
xDec#63#1 1 54 51 92 1
+ 2
+ ConvertDecode1
xDec#63#2 1 54 69 92 1
+ 2
+ ConvertDecode1
xDec#63#3 1 54 85 92 1
+ 2
+ ConvertDecode1
xDec#63#4 1 54 64 92 1
+ 2
+ ConvertDecode1
xDec#63#5 1 54 101 92 1
+ 2
+ ConvertDecode1
xDec#63#6 1 92 54 127 1
+ 2
+ ConvertDecode0
xDec#62#0 1 122 26 39 1
+ 2
+ ConvertDecode1
xDec#62#1 1 39 122 51 1
+ 2
+ ConvertDecode0
xDec#62#2 1 122 69 39 1
+ 2
+ ConvertDecode1
xDec#62#3 1 122 85 39 1
+ 2
+ ConvertDecode1
xDec#62#4 1 122 64 39 1
+ 2
+ ConvertDecode1
xDec#62#5 1 122 101 39 1
+ 2
+ ConvertDecode1
xDec#62#6 1 39 122 127 1
+ 2
+ ConvertDecode0
xDec#61#0 1 135 84 26 1
+ 2
+ ConvertDecode0
xDec#61#1 1 135 84 51 1
+ 2
+ ConvertDecode0
xDec#61#2 1 84 69 135 1
+ 2
+ ConvertDecode1
xDec#61#3 1 84 85 135 1
+ 2
+ ConvertDecode1
xDec#61#4 1 84 64 135 1
+ 2
+ ConvertDecode1
xDec#61#5 1 84 101 135 1
+ 2
+ ConvertDecode1
xDec#61#6 1 135 84 127 1
+ 2
+ ConvertDecode0
xDec#60#0 1 83 26 119 1
+ 2
+ ConvertDecode1
xDec#60#1 1 83 51 119 1
+ 2
+ ConvertDecode1
xDec#60#2 1 119 83 69 1
+ 2
+ ConvertDecode0
xDec#60#3 1 83 85 119 1
+ 2
+ ConvertDecode1
xDec#60#4 1 83 64 119 1
+ 2
+ ConvertDecode1
xDec#60#5 1 83 101 119 1
+ 2
+ ConvertDecode1
xDec#60#6 1 119 83 127 1
+ 2
+ ConvertDecode0
xDec#59#0 1 55 20 26 1
+ 2
+ ConvertDecode0
xDec#59#1 1 20 51 55 1
+ 2
+ ConvertDecode1
xDec#59#2 1 55 20 69 1
+ 2
+ ConvertDecode0
xDec#59#3 1 20 85 55 1
+ 2
+ ConvertDecode1
xDec#59#4 1 20 64 55 1
+ 2
+ ConvertDecode1
xDec#59#5 1 20 101 55 1
+ 2
+ ConvertDecode1
xDec#59#6 1 55 20 127 1
+ 2
+ ConvertDecode0
xDec#58#0 1 132 26 13 1
+ 2
+ ConvertDecode1
xDec#58#1 1 13 132 51 1
+ 2
+ ConvertDecode0
xDec#58#2 1 13 132 69 1
+ 2
+ ConvertDecode0
xDec#58#3 1 132 85 13 1
+ 2
+ ConvertDecode1
xDec#58#4 1 132 64 13 1
+ 2
+ ConvertDecode1
xDec#58#5 1 132 101 13 1
+ 2
+ ConvertDecode1
xDec#58#6 1 13 132 127 1
+ 2
+ ConvertDecode0
xDec#57#0 1 111 103 26 1
+ 2
+ ConvertDecode0
xDec#57#1 1 111 103 51 1
+ 2
+ ConvertDecode0
xDec#57#2 1 111 103 69 1
+ 2
+ ConvertDecode0
xDec#57#3 1 103 85 111 1
+ 2
+ ConvertDecode1
xDec#57#4 1 103 64 111 1
+ 2
+ ConvertDecode1
xDec#57#5 1 103 101 111 1
+ 2
+ ConvertDecode1
xDec#57#6 1 111 103 127 1
+ 2
+ ConvertDecode0
xDec#56#0 1 38 26 104 1
+ 2
+ ConvertDecode1
xDec#56#1 1 38 51 104 1
+ 2
+ ConvertDecode1
xDec#56#2 1 38 69 104 1
+ 2
+ ConvertDecode1
xDec#56#3 1 104 38 85 1
+ 2
+ ConvertDecode0
xDec#56#4 1 38 64 104 1
+ 2
+ ConvertDecode1
xDec#56#5 1 38 101 104 1
+ 2
+ ConvertDecode1
xDec#56#6 1 104 38 127 1
+ 2
+ ConvertDecode0
xDec#55#0 1 58 140 26 1
+ 2
+ ConvertDecode0
xDec#55#1 1 140 51 58 1
+ 2
+ ConvertDecode1
xDec#55#2 1 140 69 58 1
+ 2
+ ConvertDecode1
xDec#55#3 1 58 140 85 1
+ 2
+ ConvertDecode0
xDec#55#4 1 140 64 58 1
+ 2
+ ConvertDecode1
xDec#55#5 1 140 101 58 1
+ 2
+ ConvertDecode1
xDec#55#6 1 58 140 127 1
+ 2
+ ConvertDecode0
xDec#54#0 1 79 26 139 1
+ 2
+ ConvertDecode1
xDec#54#1 1 139 79 51 1
+ 2
+ ConvertDecode0
xDec#54#2 1 79 69 139 1
+ 2
+ ConvertDecode1
xDec#54#3 1 139 79 85 1
+ 2
+ ConvertDecode0
xDec#54#4 1 79 64 139 1
+ 2
+ ConvertDecode1
xDec#54#5 1 79 101 139 1
+ 2
+ ConvertDecode1
xDec#54#6 1 139 79 127 1
+ 2
+ ConvertDecode0
xDec#53#0 1 81 29 26 1
+ 2
+ ConvertDecode0
xDec#53#1 1 81 29 51 1
+ 2
+ ConvertDecode0
xDec#53#2 1 29 69 81 1
+ 2
+ ConvertDecode1
xDec#53#3 1 81 29 85 1
+ 2
+ ConvertDecode0
xDec#53#4 1 29 64 81 1
+ 2
+ ConvertDecode1
xDec#53#5 1 29 101 81 1
+ 2
+ ConvertDecode1
xDec#53#6 1 81 29 127 1
+ 2
+ ConvertDecode0
xDec#52#0 1 18 26 71 1
+ 2
+ ConvertDecode1
xDec#52#1 1 18 51 71 1
+ 2
+ ConvertDecode1
xDec#52#2 1 71 18 69 1
+ 2
+ ConvertDecode0
xDec#52#3 1 71 18 85 1
+ 2
+ ConvertDecode0
xDec#52#4 1 18 64 71 1
+ 2
+ ConvertDecode1
xDec#52#5 1 18 101 71 1
+ 2
+ ConvertDecode1
xDec#52#6 1 71 18 127 1
+ 2
+ ConvertDecode0
xDec#51#0 1 30 67 26 1
+ 2
+ ConvertDecode0
xDec#51#1 1 67 51 30 1
+ 2
+ ConvertDecode1
xDec#51#2 1 30 67 69 1
+ 2
+ ConvertDecode0
xDec#51#3 1 30 67 85 1
+ 2
+ ConvertDecode0
xDec#51#4 1 67 64 30 1
+ 2
+ ConvertDecode1
xDec#51#5 1 67 101 30 1
+ 2
+ ConvertDecode1
xDec#51#6 1 30 67 127 1
+ 2
+ ConvertDecode0
xDec#50#0 1 100 26 126 1
+ 2
+ ConvertDecode1
xDec#50#1 1 126 100 51 1
+ 2
+ ConvertDecode0
xDec#50#2 1 126 100 69 1
+ 2
+ ConvertDecode0
xDec#50#3 1 126 100 85 1
+ 2
+ ConvertDecode0
xDec#50#4 1 100 64 126 1
+ 2
+ ConvertDecode1
xDec#50#5 1 100 101 126 1
+ 2
+ ConvertDecode1
xDec#50#6 1 126 100 127 1
+ 2
+ ConvertDecode0
xDec#49#0 1 28 53 26 1
+ 2
+ ConvertDecode0
xDec#49#1 1 28 53 51 1
+ 2
+ ConvertDecode0
xDec#49#2 1 28 53 69 1
+ 2
+ ConvertDecode0
xDec#49#3 1 28 53 85 1
+ 2
+ ConvertDecode0
xDec#49#4 1 53 64 28 1
+ 2
+ ConvertDecode1
xDec#49#5 1 53 101 28 1
+ 2
+ ConvertDecode1
xDec#49#6 1 28 53 127 1
+ 2
+ ConvertDecode0
xDec#48#0 1 137 26 16 1
+ 2
+ ConvertDecode1
xDec#48#1 1 137 51 16 1
+ 2
+ ConvertDecode1
xDec#48#2 1 137 69 16 1
+ 2
+ ConvertDecode1
xDec#48#3 1 137 85 16 1
+ 2
+ ConvertDecode1
xDec#48#4 1 16 137 64 1
+ 2
+ ConvertDecode0
xDec#48#5 1 137 101 16 1
+ 2
+ ConvertDecode1
xDec#48#6 1 16 137 127 1
+ 2
+ ConvertDecode0
xDec#47#0 1 97 123 26 1
+ 2
+ ConvertDecode0
xDec#47#1 1 123 51 97 1
+ 2
+ ConvertDecode1
xDec#47#2 1 123 69 97 1
+ 2
+ ConvertDecode1
xDec#47#3 1 123 85 97 1
+ 2
+ ConvertDecode1
xDec#47#4 1 97 123 64 1
+ 2
+ ConvertDecode0
xDec#47#5 1 123 101 97 1
+ 2
+ ConvertDecode1
xDec#47#6 1 97 123 127 1
+ 2
+ ConvertDecode0
xDec#46#0 1 14 26 90 1
+ 2
+ ConvertDecode1
xDec#46#1 1 90 14 51 1
+ 2
+ ConvertDecode0
xDec#46#2 1 14 69 90 1
+ 2
+ ConvertDecode1
xDec#46#3 1 14 85 90 1
+ 2
+ ConvertDecode1
xDec#46#4 1 90 14 64 1
+ 2
+ ConvertDecode0
xDec#46#5 1 14 101 90 1
+ 2
+ ConvertDecode1
xDec#46#6 1 90 14 127 1
+ 2
+ ConvertDecode0
xDec#45#0 1 93 15 26 1
+ 2
+ ConvertDecode0
xDec#45#1 1 93 15 51 1
+ 2
+ ConvertDecode0
xDec#45#2 1 15 69 93 1
+ 2
+ ConvertDecode1
xDec#45#3 1 15 85 93 1
+ 2
+ ConvertDecode1
xDec#45#4 1 93 15 64 1
+ 2
+ ConvertDecode0
xDec#45#5 1 15 101 93 1
+ 2
+ ConvertDecode1
xDec#45#6 1 93 15 127 1
+ 2
+ ConvertDecode0
xDec#44#0 1 61 26 40 1
+ 2
+ ConvertDecode1
xDec#44#1 1 61 51 40 1
+ 2
+ ConvertDecode1
xDec#44#2 1 40 61 69 1
+ 2
+ ConvertDecode0
xDec#44#3 1 61 85 40 1
+ 2
+ ConvertDecode1
xDec#44#4 1 40 61 64 1
+ 2
+ ConvertDecode0
xDec#44#5 1 61 101 40 1
+ 2
+ ConvertDecode1
xDec#44#6 1 40 61 127 1
+ 2
+ ConvertDecode0
xDec#43#0 1 62 98 26 1
+ 2
+ ConvertDecode0
xDec#43#1 1 98 51 62 1
+ 2
+ ConvertDecode1
xDec#43#2 1 62 98 69 1
+ 2
+ ConvertDecode0
xDec#43#3 1 98 85 62 1
+ 2
+ ConvertDecode1
xDec#43#4 1 62 98 64 1
+ 2
+ ConvertDecode0
xDec#43#5 1 98 101 62 1
+ 2
+ ConvertDecode1
xDec#43#6 1 62 98 127 1
+ 2
+ ConvertDecode0
xDec#42#0 1 52 26 50 1
+ 2
+ ConvertDecode1
xDec#42#1 1 50 52 51 1
+ 2
+ ConvertDecode0
xDec#42#2 1 50 52 69 1
+ 2
+ ConvertDecode0
xDec#42#3 1 52 85 50 1
+ 2
+ ConvertDecode1
xDec#42#4 1 50 52 64 1
+ 2
+ ConvertDecode0
xDec#42#5 1 52 101 50 1
+ 2
+ ConvertDecode1
xDec#42#6 1 50 52 127 1
+ 2
+ ConvertDecode0
xDec#41#0 1 80 47 26 1
+ 2
+ ConvertDecode0
xDec#41#1 1 80 47 51 1
+ 2
+ ConvertDecode0
xDec#41#2 1 80 47 69 1
+ 2
+ ConvertDecode0
xDec#41#3 1 47 85 80 1
+ 2
+ ConvertDecode1
xDec#41#4 1 80 47 64 1
+ 2
+ ConvertDecode0
xDec#41#5 1 47 101 80 1
+ 2
+ ConvertDecode1
xDec#41#6 1 80 47 127 1
+ 2
+ ConvertDecode0
xDec#40#0 1 112 26 17 1
+ 2
+ ConvertDecode1
xDec#40#1 1 112 51 17 1
+ 2
+ ConvertDecode1
xDec#40#2 1 112 69 17 1
+ 2
+ ConvertDecode1
xDec#40#3 1 17 112 85 1
+ 2
+ ConvertDecode0
xDec#40#4 1 17 112 64 1
+ 2
+ ConvertDecode0
xDec#40#5 1 112 101 17 1
+ 2
+ ConvertDecode1
xDec#40#6 1 17 112 127 1
+ 2
+ ConvertDecode0
xDec#39#0 1 133 78 26 1
+ 2
+ ConvertDecode0
xDec#39#1 1 78 51 133 1
+ 2
+ ConvertDecode1
xDec#39#2 1 78 69 133 1
+ 2
+ ConvertDecode1
xDec#39#3 1 133 78 85 1
+ 2
+ ConvertDecode0
xDec#39#4 1 133 78 64 1
+ 2
+ ConvertDecode0
xDec#39#5 1 78 101 133 1
+ 2
+ ConvertDecode1
xDec#39#6 1 133 78 127 1
+ 2
+ ConvertDecode0
xDec#38#0 1 12 26 107 1
+ 2
+ ConvertDecode1
xDec#38#1 1 107 12 51 1
+ 2
+ ConvertDecode0
xDec#38#2 1 12 69 107 1
+ 2
+ ConvertDecode1
xDec#38#3 1 107 12 85 1
+ 2
+ ConvertDecode0
xDec#38#4 1 107 12 64 1
+ 2
+ ConvertDecode0
xDec#38#5 1 12 101 107 1
+ 2
+ ConvertDecode1
xDec#38#6 1 107 12 127 1
+ 2
+ ConvertDecode0
xDec#37#0 1 60 109 26 1
+ 2
+ ConvertDecode0
xDec#37#1 1 60 109 51 1
+ 2
+ ConvertDecode0
xDec#37#2 1 109 69 60 1
+ 2
+ ConvertDecode1
xDec#37#3 1 60 109 85 1
+ 2
+ ConvertDecode0
xDec#37#4 1 60 109 64 1
+ 2
+ ConvertDecode0
xDec#37#5 1 109 101 60 1
+ 2
+ ConvertDecode1
xDec#37#6 1 60 109 127 1
+ 2
+ ConvertDecode0
xDec#36#0 1 96 26 77 1
+ 2
+ ConvertDecode1
xDec#36#1 1 96 51 77 1
+ 2
+ ConvertDecode1
xDec#36#2 1 77 96 69 1
+ 2
+ ConvertDecode0
xDec#36#3 1 77 96 85 1
+ 2
+ ConvertDecode0
xDec#36#4 1 77 96 64 1
+ 2
+ ConvertDecode0
xDec#36#5 1 96 101 77 1
+ 2
+ ConvertDecode1
xDec#36#6 1 77 96 127 1
+ 2
+ ConvertDecode0
xDec#35#0 1 125 49 26 1
+ 2
+ ConvertDecode0
xDec#35#1 1 49 51 125 1
+ 2
+ ConvertDecode1
xDec#35#2 1 125 49 69 1
+ 2
+ ConvertDecode0
xDec#35#3 1 125 49 85 1
+ 2
+ ConvertDecode0
xDec#35#4 1 125 49 64 1
+ 2
+ ConvertDecode0
xDec#35#5 1 49 101 125 1
+ 2
+ ConvertDecode1
xDec#35#6 1 125 49 127 1
+ 2
+ ConvertDecode0
xDec#34#0 1 35 26 87 1
+ 2
+ ConvertDecode1
xDec#34#1 1 87 35 51 1
+ 2
+ ConvertDecode0
xDec#34#2 1 87 35 69 1
+ 2
+ ConvertDecode0
xDec#34#3 1 87 35 85 1
+ 2
+ ConvertDecode0
xDec#34#4 1 87 35 64 1
+ 2
+ ConvertDecode0
xDec#34#5 1 35 101 87 1
+ 2
+ ConvertDecode1
xDec#34#6 1 87 35 127 1
+ 2
+ ConvertDecode0
xDec#33#0 1 33 121 26 1
+ 2
+ ConvertDecode0
xDec#33#1 1 33 121 51 1
+ 2
+ ConvertDecode0
xDec#33#2 1 33 121 69 1
+ 2
+ ConvertDecode0
xDec#33#3 1 33 121 85 1
+ 2
+ ConvertDecode0
xDec#33#4 1 33 121 64 1
+ 2
+ ConvertDecode0
xDec#33#5 1 121 101 33 1
+ 2
+ ConvertDecode1
xDec#33#6 1 33 121 127 1
+ 2
+ ConvertDecode0
xDec#32#0 1 73 26 23 1
+ 2
+ ConvertDecode1
xDec#32#1 1 73 51 23 1
+ 2
+ ConvertDecode1
xDec#32#2 1 73 69 23 1
+ 2
+ ConvertDecode1
xDec#32#3 1 73 85 23 1
+ 2
+ ConvertDecode1
xDec#32#4 1 73 64 23 1
+ 2
+ ConvertDecode1
xDec#32#5 1 23 73 101 1
+ 2
+ ConvertDecode0
xDec#32#6 1 23 73 127 1
+ 2
+ ConvertDecode0
xDec#31#0 1 106 11 26 1
+ 2
+ ConvertDecode0
xDec#31#1 1 11 51 106 1
+ 2
+ ConvertDecode1
xDec#31#2 1 11 69 106 1
+ 2
+ ConvertDecode1
xDec#31#3 1 11 85 106 1
+ 2
+ ConvertDecode1
xDec#31#4 1 11 64 106 1
+ 2
+ ConvertDecode1
xDec#31#5 1 106 11 101 1
+ 2
+ ConvertDecode0
xDec#31#6 1 106 11 127 1
+ 2
+ ConvertDecode0
xDec#30#0 1 102 26 68 1
+ 2
+ ConvertDecode1
xDec#30#1 1 68 102 51 1
+ 2
+ ConvertDecode0
xDec#30#2 1 102 69 68 1
+ 2
+ ConvertDecode1
xDec#30#3 1 102 85 68 1
+ 2
+ ConvertDecode1
xDec#30#4 1 102 64 68 1
+ 2
+ ConvertDecode1
xDec#30#5 1 68 102 101 1
+ 2
+ ConvertDecode0
xDec#30#6 1 68 102 127 1
+ 2
+ ConvertDecode0
xDec#29#0 1 3 63 26 1
+ 2
+ ConvertDecode0
xDec#29#1 1 3 63 51 1
+ 2
+ ConvertDecode0
xDec#29#2 1 63 69 3 1
+ 2
+ ConvertDecode1
xDec#29#3 1 63 85 3 1
+ 2
+ ConvertDecode1
xDec#29#4 1 63 64 3 1
+ 2
+ ConvertDecode1
xDec#29#5 1 3 63 101 1
+ 2
+ ConvertDecode0
xDec#29#6 1 3 63 127 1
+ 2
+ ConvertDecode0
xDec#28#0 1 48 26 129 1
+ 2
+ ConvertDecode1
xDec#28#1 1 48 51 129 1
+ 2
+ ConvertDecode1
xDec#28#2 1 129 48 69 1
+ 2
+ ConvertDecode0
xDec#28#3 1 48 85 129 1
+ 2
+ ConvertDecode1
xDec#28#4 1 48 64 129 1
+ 2
+ ConvertDecode1
xDec#28#5 1 129 48 101 1
+ 2
+ ConvertDecode0
xDec#28#6 1 129 48 127 1
+ 2
+ ConvertDecode0
xDec#27#0 1 65 91 26 1
+ 2
+ ConvertDecode0
xDec#27#1 1 91 51 65 1
+ 2
+ ConvertDecode1
xDec#27#2 1 65 91 69 1
+ 2
+ ConvertDecode0
xDec#27#3 1 91 85 65 1
+ 2
+ ConvertDecode1
xDec#27#4 1 91 64 65 1
+ 2
+ ConvertDecode1
xDec#27#5 1 65 91 101 1
+ 2
+ ConvertDecode0
xDec#27#6 1 65 91 127 1
+ 2
+ ConvertDecode0
xDec#26#0 1 120 26 46 1
+ 2
+ ConvertDecode1
xDec#26#1 1 46 120 51 1
+ 2
+ ConvertDecode0
xDec#26#2 1 46 120 69 1
+ 2
+ ConvertDecode0
xDec#26#3 1 120 85 46 1
+ 2
+ ConvertDecode1
xDec#26#4 1 120 64 46 1
+ 2
+ ConvertDecode1
xDec#26#5 1 46 120 101 1
+ 2
+ ConvertDecode0
xDec#26#6 1 46 120 127 1
+ 2
+ ConvertDecode0
xDec#25#0 1 124 76 26 1
+ 2
+ ConvertDecode0
xDec#25#1 1 124 76 51 1
+ 2
+ ConvertDecode0
xDec#25#2 1 124 76 69 1
+ 2
+ ConvertDecode0
xDec#25#3 1 76 85 124 1
+ 2
+ ConvertDecode1
xDec#25#4 1 76 64 124 1
+ 2
+ ConvertDecode1
xDec#25#5 1 124 76 101 1
+ 2
+ ConvertDecode0
xDec#25#6 1 124 76 127 1
+ 2
+ ConvertDecode0
xDec#24#0 1 7 26 114 1
+ 2
+ ConvertDecode1
xDec#24#1 1 7 51 114 1
+ 2
+ ConvertDecode1
xDec#24#2 1 7 69 114 1
+ 2
+ ConvertDecode1
xDec#24#3 1 114 7 85 1
+ 2
+ ConvertDecode0
xDec#24#4 1 7 64 114 1
+ 2
+ ConvertDecode1
xDec#24#5 1 114 7 101 1
+ 2
+ ConvertDecode0
xDec#24#6 1 114 7 127 1
+ 2
+ ConvertDecode0
xDec#23#0 1 5 131 26 1
+ 2
+ ConvertDecode0
xDec#23#1 1 131 51 5 1
+ 2
+ ConvertDecode1
xDec#23#2 1 131 69 5 1
+ 2
+ ConvertDecode1
xDec#23#3 1 5 131 85 1
+ 2
+ ConvertDecode0
xDec#23#4 1 131 64 5 1
+ 2
+ ConvertDecode1
xDec#23#5 1 5 131 101 1
+ 2
+ ConvertDecode0
xDec#23#6 1 5 131 127 1
+ 2
+ ConvertDecode0
xDec#22#0 1 56 26 21 1
+ 2
+ ConvertDecode1
xDec#22#1 1 21 56 51 1
+ 2
+ ConvertDecode0
xDec#22#2 1 56 69 21 1
+ 2
+ ConvertDecode1
xDec#22#3 1 21 56 85 1
+ 2
+ ConvertDecode0
xDec#22#4 1 56 64 21 1
+ 2
+ ConvertDecode1
xDec#22#5 1 21 56 101 1
+ 2
+ ConvertDecode0
xDec#22#6 1 21 56 127 1
+ 2
+ ConvertDecode0
xDec#21#0 1 128 45 26 1
+ 2
+ ConvertDecode0
xDec#21#1 1 128 45 51 1
+ 2
+ ConvertDecode0
xDec#21#2 1 45 69 128 1
+ 2
+ ConvertDecode1
xDec#21#3 1 128 45 85 1
+ 2
+ ConvertDecode0
xDec#21#4 1 45 64 128 1
+ 2
+ ConvertDecode1
xDec#21#5 1 128 45 101 1
+ 2
+ ConvertDecode0
xDec#21#6 1 128 45 127 1
+ 2
+ ConvertDecode0
xDec#20#0 1 27 26 108 1
+ 2
+ ConvertDecode1
xDec#20#1 1 27 51 108 1
+ 2
+ ConvertDecode1
xDec#20#2 1 108 27 69 1
+ 2
+ ConvertDecode0
xDec#20#3 1 108 27 85 1
+ 2
+ ConvertDecode0
xDec#20#4 1 27 64 108 1
+ 2
+ ConvertDecode1
xDec#20#5 1 108 27 101 1
+ 2
+ ConvertDecode0
xDec#20#6 1 108 27 127 1
+ 2
+ ConvertDecode0
xDec#19#0 1 24 117 26 1
+ 2
+ ConvertDecode0
xDec#19#1 1 117 51 24 1
+ 2
+ ConvertDecode1
xDec#19#2 1 24 117 69 1
+ 2
+ ConvertDecode0
xDec#19#3 1 24 117 85 1
+ 2
+ ConvertDecode0
xDec#19#4 1 117 64 24 1
+ 2
+ ConvertDecode1
xDec#19#5 1 24 117 101 1
+ 2
+ ConvertDecode0
xDec#19#6 1 24 117 127 1
+ 2
+ ConvertDecode0
xDec#18#0 1 66 26 9 1
+ 2
+ ConvertDecode1
xDec#18#1 1 9 66 51 1
+ 2
+ ConvertDecode0
xDec#18#2 1 9 66 69 1
+ 2
+ ConvertDecode0
xDec#18#3 1 9 66 85 1
+ 2
+ ConvertDecode0
xDec#18#4 1 66 64 9 1
+ 2
+ ConvertDecode1
xDec#18#5 1 9 66 101 1
+ 2
+ ConvertDecode0
xDec#18#6 1 9 66 127 1
+ 2
+ ConvertDecode0
xDec#17#0 1 95 6 26 1
+ 2
+ ConvertDecode0
xDec#17#1 1 95 6 51 1
+ 2
+ ConvertDecode0
xDec#17#2 1 95 6 69 1
+ 2
+ ConvertDecode0
xDec#17#3 1 95 6 85 1
+ 2
+ ConvertDecode0
xDec#17#4 1 6 64 95 1
+ 2
+ ConvertDecode1
xDec#17#5 1 95 6 101 1
+ 2
+ ConvertDecode0
xDec#17#6 1 95 6 127 1
+ 2
+ ConvertDecode0
xDec#16#0 1 94 26 88 1
+ 2
+ ConvertDecode1
xDec#16#1 1 94 51 88 1
+ 2
+ ConvertDecode1
xDec#16#2 1 94 69 88 1
+ 2
+ ConvertDecode1
xDec#16#3 1 94 85 88 1
+ 2
+ ConvertDecode1
xDec#16#4 1 88 94 64 1
+ 2
+ ConvertDecode0
xDec#16#5 1 88 94 101 1
+ 2
+ ConvertDecode0
xDec#16#6 1 88 94 127 1
+ 2
+ ConvertDecode0
xDec#15#0 1 34 57 26 1
+ 2
+ ConvertDecode0
xDec#15#1 1 57 51 34 1
+ 2
+ ConvertDecode1
xDec#15#2 1 57 69 34 1
+ 2
+ ConvertDecode1
xDec#15#3 1 57 85 34 1
+ 2
+ ConvertDecode1
xDec#15#4 1 34 57 64 1
+ 2
+ ConvertDecode0
xDec#15#5 1 34 57 101 1
+ 2
+ ConvertDecode0
xDec#15#6 1 34 57 127 1
+ 2
+ ConvertDecode0
xDec#14#0 1 42 26 134 1
+ 2
+ ConvertDecode1
xDec#14#1 1 134 42 51 1
+ 2
+ ConvertDecode0
xDec#14#2 1 42 69 134 1
+ 2
+ ConvertDecode1
xDec#14#3 1 42 85 134 1
+ 2
+ ConvertDecode1
xDec#14#4 1 134 42 64 1
+ 2
+ ConvertDecode0
xDec#14#5 1 134 42 101 1
+ 2
+ ConvertDecode0
xDec#14#6 1 134 42 127 1
+ 2
+ ConvertDecode0
xDec#13#0 1 59 86 26 1
+ 2
+ ConvertDecode0
xDec#13#1 1 59 86 51 1
+ 2
+ ConvertDecode0
xDec#13#2 1 86 69 59 1
+ 2
+ ConvertDecode1
xDec#13#3 1 86 85 59 1
+ 2
+ ConvertDecode1
xDec#13#4 1 59 86 64 1
+ 2
+ ConvertDecode0
xDec#13#5 1 59 86 101 1
+ 2
+ ConvertDecode0
xDec#13#6 1 59 86 127 1
+ 2
+ ConvertDecode0
xDec#12#0 1 115 26 44 1
+ 2
+ ConvertDecode1
xDec#12#1 1 115 51 44 1
+ 2
+ ConvertDecode1
xDec#12#2 1 44 115 69 1
+ 2
+ ConvertDecode0
xDec#12#3 1 115 85 44 1
+ 2
+ ConvertDecode1
xDec#12#4 1 44 115 64 1
+ 2
+ ConvertDecode0
xDec#12#5 1 44 115 101 1
+ 2
+ ConvertDecode0
xDec#12#6 1 44 115 127 1
+ 2
+ ConvertDecode0
xDec#11#0 1 4 72 26 1
+ 2
+ ConvertDecode0
xDec#11#1 1 72 51 4 1
+ 2
+ ConvertDecode1
xDec#11#2 1 4 72 69 1
+ 2
+ ConvertDecode0
xDec#11#3 1 72 85 4 1
+ 2
+ ConvertDecode1
xDec#11#4 1 4 72 64 1
+ 2
+ ConvertDecode0
xDec#11#5 1 4 72 101 1
+ 2
+ ConvertDecode0
xDec#11#6 1 4 72 127 1
+ 2
+ ConvertDecode0
xDec#10#0 1 138 26 36 1
+ 2
+ ConvertDecode1
xDec#10#1 1 36 138 51 1
+ 2
+ ConvertDecode0
xDec#10#2 1 36 138 69 1
+ 2
+ ConvertDecode0
xDec#10#3 1 138 85 36 1
+ 2
+ ConvertDecode1
xDec#10#4 1 36 138 64 1
+ 2
+ ConvertDecode0
xDec#10#5 1 36 138 101 1
+ 2
+ ConvertDecode0
xDec#10#6 1 36 138 127 1
+ 2
+ ConvertDecode0
xDec#9#0 1 136 118 26 1
+ 2
+ ConvertDecode0
xDec#9#1 1 136 118 51 1
+ 2
+ ConvertDecode0
xDec#9#2 1 136 118 69 1
+ 2
+ ConvertDecode0
xDec#9#3 1 118 85 136 1
+ 2
+ ConvertDecode1
xDec#9#4 1 136 118 64 1
+ 2
+ ConvertDecode0
xDec#9#5 1 136 118 101 1
+ 2
+ ConvertDecode0
xDec#9#6 1 136 118 127 1
+ 2
+ ConvertDecode0
xDec#8#0 1 41 26 113 1
+ 2
+ ConvertDecode1
xDec#8#1 1 41 51 113 1
+ 2
+ ConvertDecode1
xDec#8#2 1 41 69 113 1
+ 2
+ ConvertDecode1
xDec#8#3 1 113 41 85 1
+ 2
+ ConvertDecode0
xDec#8#4 1 113 41 64 1
+ 2
+ ConvertDecode0
xDec#8#5 1 113 41 101 1
+ 2
+ ConvertDecode0
xDec#8#6 1 113 41 127 1
+ 2
+ ConvertDecode0
xDec#7#0 1 75 8 26 1
+ 2
+ ConvertDecode0
xDec#7#1 1 8 51 75 1
+ 2
+ ConvertDecode1
xDec#7#2 1 8 69 75 1
+ 2
+ ConvertDecode1
xDec#7#3 1 75 8 85 1
+ 2
+ ConvertDecode0
xDec#7#4 1 75 8 64 1
+ 2
+ ConvertDecode0
xDec#7#5 1 75 8 101 1
+ 2
+ ConvertDecode0
xDec#7#6 1 75 8 127 1
+ 2
+ ConvertDecode0
xDec#6#0 1 82 26 10 1
+ 2
+ ConvertDecode1
xDec#6#1 1 10 82 51 1
+ 2
+ ConvertDecode0
xDec#6#2 1 82 69 10 1
+ 2
+ ConvertDecode1
xDec#6#3 1 10 82 85 1
+ 2
+ ConvertDecode0
xDec#6#4 1 10 82 64 1
+ 2
+ ConvertDecode0
xDec#6#5 1 10 82 101 1
+ 2
+ ConvertDecode0
xDec#6#6 1 10 82 127 1
+ 2
+ ConvertDecode0
xDec#5#0 1 130 32 26 1
+ 2
+ ConvertDecode0
xDec#5#1 1 130 32 51 1
+ 2
+ ConvertDecode0
xDec#5#2 1 32 69 130 1
+ 2
+ ConvertDecode1
xDec#5#3 1 130 32 85 1
+ 2
+ ConvertDecode0
xDec#5#4 1 130 32 64 1
+ 2
+ ConvertDecode0
xDec#5#5 1 130 32 101 1
+ 2
+ ConvertDecode0
xDec#5#6 1 130 32 127 1
+ 2
+ ConvertDecode0
xDec#4#0 1 43 26 99 1
+ 2
+ ConvertDecode1
xDec#4#1 1 43 51 99 1
+ 2
+ ConvertDecode1
xDec#4#2 1 99 43 69 1
+ 2
+ ConvertDecode0
xDec#4#3 1 99 43 85 1
+ 2
+ ConvertDecode0
xDec#4#4 1 99 43 64 1
+ 2
+ ConvertDecode0
xDec#4#5 1 99 43 101 1
+ 2
+ ConvertDecode0
xDec#4#6 1 99 43 127 1
+ 2
+ ConvertDecode0
xDec#3#0 1 31 70 26 1
+ 2
+ ConvertDecode0
xDec#3#1 1 70 51 31 1
+ 2
+ ConvertDecode1
xDec#3#2 1 31 70 69 1
+ 2
+ ConvertDecode0
xDec#3#3 1 31 70 85 1
+ 2
+ ConvertDecode0
xDec#3#4 1 31 70 64 1
+ 2
+ ConvertDecode0
xDec#3#5 1 31 70 101 1
+ 2
+ ConvertDecode0
xDec#3#6 1 31 70 127 1
+ 2
+ ConvertDecode0
xDec#2#0 1 116 26 19 1
+ 2
+ ConvertDecode1
xDec#2#1 1 19 116 51 1
+ 2
+ ConvertDecode0
xDec#2#2 1 19 116 69 1
+ 2
+ ConvertDecode0
xDec#2#3 1 19 116 85 1
+ 2
+ ConvertDecode0
xDec#2#4 1 19 116 64 1
+ 2
+ ConvertDecode0
xDec#2#5 1 19 116 101 1
+ 2
+ ConvertDecode0
xDec#2#6 1 19 116 127 1
+ 2
+ ConvertDecode0
xDec#1#0 1 22 74 26 1
+ 2
+ ConvertDecode0
xDec#1#1 1 22 74 51 1
+ 2
+ ConvertDecode0
xDec#1#2 1 22 74 69 1
+ 2
+ ConvertDecode0
xDec#1#3 1 22 74 85 1
+ 2
+ ConvertDecode0
xDec#1#4 1 22 74 64 1
+ 2
+ ConvertDecode0
xDec#1#5 1 22 74 101 1
+ 2
+ ConvertDecode0
xDec#1#6 1 22 74 127 1
+ 2
+ ConvertDecode0
xDec#0#0 1 37 110 26 1
+ 2
+ ConvertDecode0
xDec#0#1 1 37 110 51 1
+ 2
+ ConvertDecode0
xDec#0#2 1 37 110 69 1
+ 2
+ ConvertDecode0
xDec#0#3 1 37 110 85 1
+ 2
+ ConvertDecode0
xDec#0#4 1 37 110 64 1
+ 2
+ ConvertDecode0
xDec#0#5 1 37 110 101 1
+ 2
+ ConvertDecode0
xDec#0#6 1 110 127 37 1
+ 2
+ ConvertDecode1
.ends ConvertDecode
.subckt ConDecRtg 1 2 3 4 5
+ 6 7 8 9 10 11
+ 12 13 14 15 16
c426 13 15 5.34017e-13
c427 14 15 1.06691e-12
c428 12 15 9.91344e-13
c429 11 15 5.53835e-13
c430 9 15 5.36293e-13
c431 10 15 7.45956e-13
c432 8 15 6.70388e-13
c433 7 15 5.5611e-13
c434 5 15 5.38568e-13
c435 6 15 4.25001e-13
c436 4 15 3.49432e-13
c437 3 15 5.58387e-13
c438 1 15 5.40845e-13
c439 2 15 1.04045e-13
c440 3 14 1.75e-14
c441 7 14 1.75e-14
c442 3 9 1.75e-14
c443 7 9 1.75e-14
c444 3 6 1.75e-14
c445 5 11 1.75e-14
c446 3 7 1.75e-14
c447 3 8 1.75e-14
c448 1 14 1.75e-14
c449 7 8 1.75e-14
c450 1 9 1.75e-14
c451 1 6 1.75e-14
c452 5 12 1.75e-14
c453 5 10 1.75e-14
c454 1 3 1.75e-14
c455 1 7 1.75e-14
c456 1 8 1.75e-14
c457 9 13 1.75e-14
c458 11 14 1.75e-14
c459 3 13 1.75e-14
c460 9 11 1.75e-14
c461 7 13 1.75e-14
c462 3 11 1.75e-14
c463 7 11 1.75e-14
c464 9 12 1.75e-14
c465 1 13 1.75e-14
c466 5 14 1.75e-14
c467 3 12 1.75e-14
c468 7 12 1.75e-14
c469 5 9 1.75e-14
c470 1 11 1.75e-14
c471 3 10 1.75e-14
c472 7 10 1.75e-14
c473 3 5 1.75e-14
c474 5 7 1.75e-14
c475 5 8 1.75e-14
c476 1 12 1.75e-14
c477 11 13 1.75e-14
c478 1 10 1.75e-14
c479 3 4 1.75e-14
c480 1 5 1.75e-14
c481 1 4 1.75e-14
c482 9 14 1.75e-14
c483 11 12 1.75e-14
c484 5 13 1.75e-14
.ends ConDecRtg
.subckt AtoDRtgE 1 2 3 4 5
+ 6 7 8 9 10 11
+ 12 13 14
c485 8 9 7.66022e-11
c486 7 9 2.27177e-12
c487 6 9 2.27177e-12
c488 5 9 2.27177e-12
c489 4 9 2.27177e-12
c490 3 9 2.27177e-12
c491 2 9 2.27177e-12
c492 1 9 2.27177e-12
c493 9 13 4.90118e-12
c494 9 12 4.88995e-12
c495 9 11 4.87871e-12
c496 9 10 4.87871e-12
c497 8 11 4.2e-13
c498 2 8 1.68e-12
c499 5 11 4.9e-14
c500 11 13 4.2e-14
c501 11 14 1.2e-13
c502 3 8 1.68e-12
c503 2 13 4.9e-14
c504 2 14 1.4e-13
c505 3 13 4.9e-14
c506 3 14 1.4e-13
c507 2 11 4.9e-14
c508 3 11 4.9e-14
c509 8 10 4.2e-13
c510 5 10 4.9e-14
c511 6 12 4.9e-14
c512 10 14 2.4e-13
c513 10 13 4.2e-14
c514 10 11 4.2e-14
c515 2 10 4.9e-14
c516 3 10 4.9e-14
c517 7 12 4.9e-14
c518 4 12 4.9e-14
c519 1 12 4.9e-14
c520 6 8 1.68e-12
c521 6 13 4.9e-14
c522 6 14 1.4e-13
c523 6 11 4.9e-14
c524 7 8 1.68e-12
c525 4 8 1.68e-12
c526 7 14 1.4e-13
c527 7 13 4.9e-14
c528 4 13 4.9e-14
c529 4 14 1.4e-13
c530 1 8 1.68e-12
c531 7 11 4.9e-14
c532 6 10 4.9e-14
c533 4 11 4.9e-14
c534 1 14 1.4e-13
c535 1 13 4.9e-14
c536 1 11 4.9e-14
c537 8 12 4.2e-13
c538 5 12 4.9e-14
c539 7 10 4.9e-14
c540 12 14 1.2e-13
c541 12 13 4.2e-14
c542 4 10 4.9e-14
c543 11 12 4.2e-14
c544 2 12 4.9e-14
c545 1 10 4.9e-14
c546 3 12 4.9e-14
c547 10 12 4.2e-14
c548 5 8 1.68e-12
c549 8 14 1.2e-12
c550 8 13 4.2e-13
c551 5 14 1.4e-13
c552 5 13 4.9e-14
c553 13 14 1.2e-13
.ends AtoDRtgE
xz2xCMP#0#0 0 1 3 4 5
+ 6 7 8 9 10 11 z2xCMP
xz2xCMP#0#1 0 1 16 17 18
+ 19 7 9 20 10 11 z2xCMP
xz2xCMP#0#2 0 1 25 26 27
+ 28 7 20 29 10 11 z2xCMP
xz2xCMP#0#3 0 1 34 35 36
+ 37 7 29 38 10 11 z2xCMP
xz2xCMP#0#4 0 1 43 44 45
+ 46 7 38 47 10 11 z2xCMP
xz2xCMP#0#5 0 1 52 53 54
+ 55 7 47 56 10 11 z2xCMP
xz2xCMP#0#6 0 1 61 62 63
+ 64 7 56 65 10 11 z2xCMP
xz2xCMP#0#7 0 1 70 71 72
+ 73 7 65 74 10 11 z2xCMP
xz2xCMP#0#8 0 1 79 80 81
+ 82 7 74 83 10 11 z2xCMP
xz2xCMP#0#9 0 1 88 89 90
+ 91 7 83 92 10 11 z2xCMP
xz2xCMP#0#10 0 1 97 98 99
+ 100 7 92 101 10 11 z2xCMP
xz2xCMP#0#11 0 1 106 107 108
+ 109 7 101 110 10 11 z2xCMP
xz2xCMP#0#12 0 1 115 116 117
+ 118 7 110 119 10 11 z2xCMP
xz2xCMP#0#13 0 1 124 125 126
+ 127 7 119 128 10 11 z2xCMP
xz2xCMP#0#14 0 1 133 134 135
+ 136 7 128 137 10 11 z2xCMP
xz2xCMP#0#15 0 1 142 143 144
+ 145 7 137 146 10 11 z2xCMP
xz2xCMP#0#16 0 1 151 152 153
+ 154 7 146 155 10 11 z2xCMP
xz2xCMP#0#17 0 1 160 161 162
+ 163 7 155 164 10 11 z2xCMP
xz2xCMP#0#18 0 1 169 170 171
+ 172 7 164 173 10 11 z2xCMP
xz2xCMP#0#19 0 1 178 179 180
+ 181 7 173 182 10 11 z2xCMP
xz2xCMP#0#20 0 1 187 188 189
+ 190 7 182 191 10 11 z2xCMP
xz2xCMP#0#21 0 1 196 197 198
+ 199 7 191 200 10 11 z2xCMP
xz2xCMP#0#22 0 1 205 206 207
+ 208 7 200 209 10 11 z2xCMP
xz2xCMP#0#23 0 1 214 215 216
+ 217 7 209 218 10 11 z2xCMP
xz2xCMP#0#24 0 1 223 224 225
+ 226 7 218 227 10 11 z2xCMP
xz2xCMP#0#25 0 1 232 233 234
+ 235 7 227 236 10 11 z2xCMP
xz2xCMP#0#26 0 1 241 242 243
+ 244 7 236 245 10 11 z2xCMP
xz2xCMP#0#27 0 1 250 251 252
+ 253 7 245 254 10 11 z2xCMP
xz2xCMP#0#28 0 1 259 260 261
+ 262 7 254 263 10 11 z2xCMP
xz2xCMP#0#29 0 1 268 269 270
+ 271 7 263 272 10 11 z2xCMP
xz2xCMP#0#30 0 1 277 278 279
+ 280 7 272 281 10 11 z2xCMP
xz2xCMP#0#31 0 1 286 287 288
+ 289 7 281 290 10 11 z2xCMP
xAVddRtg#0 1 0 1 AVddRtg
xCMP#0 290 10 1 7 11
+ 295 0 296 1 CMP
xFlashLatchBlnk#0 0 299 300 301 302
+ 1
+ FlashLatchBlnk
xFlashOneHot#0 0 1 214 188 107
+ 142 116 88 223 16 4
+ 151 89 224 61 35 17
+ 259 233 152 187 161 3
+ 268 115 299 196 269 124
+ 80 62 278 197 34 232
+ 206 125 160 134 241 169
+ 242 53 79 296 277 251
+ 170 179 205 286 133 287
+ 215 52 26 250 143 178
+ 106 260 71 25 97 98
+ 70 44 43 153 303 304
+ 127 305 135 279 306 109
+ 5 307 253 308 309 261
+ 310 311 235 312 198 313
+ 300 172 180 314 45 154
+ 54 19 315 28 280 316
+ 117 317 318 99 319 320
+ 243 321 322 217 323 225
+ 324 90 325 326 199 64
+ 327 73 328 329 162 136
+ 144 288 330 118 18 262
+ 301 331 270 332 244 333
+ 334 335 336 207 337 181
+ 189 338 339 163 63 340
+ 37 341 289 126 302 342
+ 100 108 252 343 226 234
+ 344 208 82 345 171 346
+ 145 347 27 348 271 349
+ 350 351 352 216 353 190
+ 72 46 354 355 356 357
+ 358 359 360 361 362 363
+ 91 36 6 364 81 365
+ 55 366 367 368 295 FlashOneHot
xz7xConvertLatch#0 0 1 299 300 301
+ 302 1085 1086 1087 1088 1089
+ 1090 1091 1092 1093 1094 1095
+ 1096 1097 1098 z7xConvertLatch
xAtoDRtgW#0 10 7 11 0 1 AtoDRtgW
xConvertDecode#0 0 1 134 53 107
+ 303 304 305 88 34 306
+ 307 268 308 309 223 187
+ 310 16 311 106 4 151
+ 89 296 1087 312 224 313
+ 233 17 314 152 71 315
+ 52 3 316 286 205 317
+ 318 319 61 320 124 321
+ 322 323 196 1090 324 325
+ 326 269 327 328 251 62
+ 170 329 197 330 1092 125
+ 331 332 142 1093 333 241
+ 334 335 336 35 337 169
+ 338 339 188 242 340 341
+ 342 1096 343 160 79 344
+ 214 345 287 206 346 80
+ 347 215 348 25 349 1097
+ 350 351 259 352 143 178
+ 97 353 354 260 355 43
+ 115 356 357 358 359 277
+ 360 361 362 363 116 161
+ 232 1098 98 133 26 364
+ 365 179 70 278 44 366
+ 367 250 368 ConvertDecode
xConDecRtg#0 1085 1087 1094 1090 1088
+ 1093 1095 1096 1089 1092 1086
+ 1097 1091 1098 0 1 ConDecRtg
xAtoDRtgE#0 1085 1094 1088 1095 1089
+ 1086 1091 1 0 299 300
+ 301 302 1 AtoDRtgE
c554 10 0 3.3696e-14
c555 1091 0 3.5e-14
c556 1086 0 3.5e-14
c557 1089 0 3.5e-14
c558 1095 0 3.5e-14
c559 1088 0 3.5e-14
c560 1094 0 3.5e-14
c561 1085 0 3.5e-14
c562 11 0 4e-14
c563 0 302 1.225e-13
c564 0 301 1.225e-13
c565 0 300 1.225e-13
c566 0 299 1.225e-13
c567 0 296 1.5625e-14
c568 0 287 1.5625e-14
c569 0 286 1.5625e-14
c570 0 278 1.5625e-14
c571 0 277 1.5625e-14
c572 0 269 1.5625e-14
c573 0 268 1.5625e-14
c574 0 260 1.5625e-14
c575 0 259 1.5625e-14
c576 0 251 1.5625e-14
c577 0 250 1.5625e-14
c578 0 242 1.5625e-14
c579 0 241 1.5625e-14
c580 0 233 1.5625e-14
c581 0 232 1.5625e-14
c582 0 224 1.5625e-14
c583 0 223 1.5625e-14
c584 0 215 1.5625e-14
c585 0 214 1.5625e-14
c586 0 206 1.5625e-14
c587 0 205 1.5625e-14
c588 0 197 1.5625e-14
c589 0 196 1.5625e-14
c590 0 188 1.5625e-14
c591 0 187 1.5625e-14
c592 0 179 1.5625e-14
c593 0 178 1.5625e-14
c594 0 170 1.5625e-14
c595 0 169 1.5625e-14
c596 0 161 1.5625e-14
c597 0 160 1.5625e-14
c598 0 152 1.5625e-14
c599 0 151 1.5625e-14
c600 0 143 1.5625e-14
c601 0 142 1.5625e-14
c602 0 134 1.5625e-14
c603 0 133 1.5625e-14
c604 0 125 1.5625e-14
c605 0 124 1.5625e-14
c606 0 116 1.5625e-14
c607 0 115 1.5625e-14
c608 0 107 1.5625e-14
c609 0 106 1.5625e-14
c610 0 98 1.5625e-14
c611 0 97 1.5625e-14
c612 0 89 1.5625e-14
c613 0 88 1.5625e-14
c614 0 80 1.5625e-14
c615 0 79 1.5625e-14
c616 0 71 1.5625e-14
c617 0 70 1.5625e-14
c618 0 62 1.5625e-14
c619 0 61 1.5625e-14
c620 0 53 1.5625e-14
c621 0 52 1.5625e-14
c622 0 44 1.5625e-14
c623 0 43 1.5625e-14
c624 0 35 1.5625e-14
c625 0 34 1.5625e-14
c626 0 26 1.5625e-14
c627 0 25 1.5625e-14
c628 0 17 1.5625e-14
c629 0 16 1.5625e-14
c630 0 4 1.5625e-14
c631 0 3 1.5625e-14
c632 7 0 1.5625e-14
c636 8 0 1e-15
VTapA0 3 0 pwl (0 0 1e-08 5 1e-07 5 1.1e-07 0 
+ 1.5e-07 10 2e-07 0 )
VVDD 1 0 5
.print TRAN v(3) v(1085) v(1094) v(1088) v(1095) v(1089) 
+v(1086) v(1091) 
.options limpts=50000 itl5=50000
.TRAN 2e-09 2e-07
.end
